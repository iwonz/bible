GEN|1|1|На початку Бог створив Небо та землю.
GEN|1|2|А земля була пуста та порожня, і темрява була над безоднею, і Дух Божий ширяв над поверхнею води.
GEN|1|3|І сказав Бог: Хай станеться світло! І сталося світло.
GEN|1|4|І побачив Бог світло, що добре воно, і Бог відділив світло від темряви.
GEN|1|5|І Бог назвав світло: День, а темряву назвав: Ніч. І був вечір, і був ранок, день перший.
GEN|1|6|І сказав Бог: Нехай станеться твердь посеред води, і нехай відділяє вона між водою й водою.
GEN|1|7|І Бог твердь учинив, і відділив воду, що під твердю вона, і воду, що над твердю вона. І сталося так.
GEN|1|8|І назвав Бог твердь Небо. І був вечір, і був ранок день другий.
GEN|1|9|І сказав Бог: Нехай збереться вода з-попід неба до місця одного, і нехай суходіл стане видний. І сталося так.
GEN|1|10|І назвав Бог суходіл: Земля, а місце зібрання води назвав: Море. І Бог побачив, що добре воно.
GEN|1|11|І сказав Бог: Нехай земля вродить траву, ярину, що насіння вона розсіває, дерево овочеве, що за родом своїм плід приносить, що в ньому насіння його на землі. І сталося так.
GEN|1|12|І земля траву видала, ярину, що насіння розсіває за родом її, і дерево, що приносить плід, що насіння його в нім за родом його. І Бог побачив, що добре воно.
GEN|1|13|І був вечір, і був ранок, день третій.
GEN|1|14|І сказав Бог: Нехай будуть світила на тверді небесній для відділення дня від ночі, і нехай вони стануть знаками, і часами умовленими, і днями, і роками.
GEN|1|15|І нехай вони стануть на тверді небесній світилами, щоб світити над землею. І сталося так.
GEN|1|16|І вчинив Бог обидва світила великі, світило велике, щоб воно керувало днем, і світило мале, щоб керувало ніччю, також зорі.
GEN|1|17|І Бог умістив їх на тверді небесній, щоб світили вони над землею,
GEN|1|18|і щоб керували днем та ніччю, і щоб відділювали світло від темряви. І Бог побачив, що це добре.
GEN|1|19|І був вечір, і був ранок, день четвертий.
GEN|1|20|І сказав Бог: Нехай вода вироїть дрібні істоти, душу живу, і птаство, що літає над землею під небесною твердю.
GEN|1|21|І створив Бог риби великі, і всяку душу живу плазуючу, що її вода вироїла за їх родом, і всяку пташину крилату за родом її. І Бог побачив, що добре воно.
GEN|1|22|І поблагословив їх Бог, кажучи: Плодіться й розмножуйтеся, і наповнюйте воду в морях, а птаство нехай розмножується на землі!
GEN|1|23|І був вечір, і був ранок, день п'ятий.
GEN|1|24|І сказав Бог: Нехай видасть земля живу душу за родом її, худобу й плазуюче, і земну звірину за родом її. І сталося так.
GEN|1|25|І вчинив Бог земну звірину за родом її, і худобу за родом її, і все земне плазуюче за родом його. І бачив Бог, що добре воно.
GEN|1|26|І сказав Бог: Створімо людину за образом Нашим, за подобою Нашою, і хай панують над морською рибою, і над птаством небесним, і над худобою, і над усею землею, і над усім плазуючим, що плазує по землі.
GEN|1|27|І Бог на Свій образ людину створив, на образ Божий її Він створив, як чоловіка та жінку створив їх.
GEN|1|28|І поблагословив їх Бог, і сказав Бог до них: Плодіться й розмножуйтеся, і наповнюйте землю, оволодійте нею, і пануйте над морськими рибами, і над птаством небесним, і над кожним плазуючим живим на землі!
GEN|1|29|І сказав Бог: Оце дав Я вам усю ярину, що розсіває насіння, що на всій землі, і кожне дерево, що на ньому плід деревний, що воно розсіває насіння, нехай буде на їжу це вам!
GEN|1|30|І земній усій звірині і всьому птаству небесному, і кожному, що плазує по землі, що душа в ньому жива, уся зелень яринна на їжу для них. І сталося так.
GEN|1|31|І побачив Бог усе, що вчинив. І ото, вельми добре воно! І був вечір, і був ранок, день шостий.
GEN|2|1|І були скінчені небо й земля, і все воїнство їхнє.
GEN|2|2|І скінчив Бог дня сьомого працю Свою, яку Він чинив. І Він відпочив у дні сьомім від усієї праці Своєї, яку був чинив.
GEN|2|3|І поблагословив Бог день сьомий, і його освятив, бо в нім відпочив Він від усієї праці Своєї, яку, чинячи, Бог був створив.
GEN|2|4|Це ось походження неба й землі, коли створено їх, у дні, як Господь Бог создав небо та землю.
GEN|2|5|І не було на землі жодної польової рослини, і жодна ярина польова не росла, бо на землю дощу Господь Бог не давав, і не було людини, щоб порати землю.
GEN|2|6|І пара з землі підіймалась, і напувала всю землю.
GEN|2|7|І створив Господь Бог людину з пороху земного. І дихання життя вдихнув у ніздрі її, і стала людина живою душею.
GEN|2|8|І насадив Господь Бог рай ув Едені на сході, і там осадив людину, що її Він створив.
GEN|2|9|І зростив Господь Бог із землі кожне дерево, принадне на вигляд і на їжу смачне, і дерево життя посеред раю, і дерево Пізнання добра і зла.
GEN|2|10|І річка з Едену виходить, щоб поїти рай. І звідти розділюється і стає чотирма початками.
GEN|2|11|Імення одному Пішон, оточує він усю землю Хавіла, де є золото.
GEN|2|12|А золото тієї землі добре; там бделій і камінь онікс.
GEN|2|13|Ім'я ж другої річки Ґіхон, вона оточує ввесь край Етіопії.
GEN|2|14|А ім'я річки третьої Тигр, вона протікає на сході Ашшуру. А річка четверта вона Ефрат.
GEN|2|15|І взяв Господь Бог людину, і в еденському раї вмістив був її, щоб порала його та його доглядала.
GEN|2|16|І наказав Господь Бог Адамові, кажучи: Із кожного дерева в Раю ти можеш їсти.
GEN|2|17|Але з дерева знання добра й зла не їж від нього, бо в день їди твоєї від нього ти напевно помреш!
GEN|2|18|І сказав Господь Бог: Не добре, щоб бути чоловіку самотнім. Створю йому поміч, подібну до нього.
GEN|2|19|І вчинив Господь Бог із землі всю польову звірину, і все птаство небесне, і до Адама привів, щоб побачити, як він їх кликатиме. А все, як покличе Адам до них, до живої душі воно ймення йому.
GEN|2|20|І назвав Адам імена всій худобі, і птаству небесному, і всій польовій звірині. Але Адамові помочі Він не знайшов, щоб подібна до нього була.
GEN|2|21|І вчинив Господь Бог, що на Адама спав міцний сон, і заснув він. І Він узяв одне з ребер його, і тілом закрив його місце.
GEN|2|22|І перетворив Господь Бог те ребро, що взяв із Адама, на жінку, і привів її до Адама.
GEN|2|23|І промовив Адам: Оце тепер вона кість від костей моїх, і тіло від тіла мого. Вона чоловіковою буде зватися, бо взята вона з чоловіка.
GEN|2|24|Покине тому чоловік свого батька та матір свою, та й пристане до жінки своєї, і стануть вони одним тілом.
GEN|2|25|І були вони нагі обоє, Адам та жінка його, і вони не соромились.
GEN|3|1|Але змій був хитріший над усю польову звірину, яку Господь Бог учинив. І сказав він до жінки: Чи Бог наказав: Не їжте з усякого дерева раю?
GEN|3|2|І відповіла жінка змієві: З плодів дерева раю ми можемо їсти,
GEN|3|3|але з плодів дерева, що в середині раю, Бог сказав: Не їжте із нього, і не доторкайтесь до нього, щоб вам не померти.
GEN|3|4|І сказав змій до жінки: Умерти не вмрете!
GEN|3|5|Бо відає Бог, що дня того, коли будете з нього ви їсти, ваші очі розкриються, і станете ви, немов Боги, знаючи добро й зло.
GEN|3|6|І побачила жінка, що дерево добре на їжу, і принадне для очей, і пожадане дерево, щоб набути знання. І взяла з його плоду, та й з'їла, і разом дала теж чоловікові своєму, і він з'їв.
GEN|3|7|І розкрилися очі в обох них, і пізнали, що нагі вони. І зшили вони фіґові листя, і зробили опаски собі.
GEN|3|8|І почули вони голос Господа Бога, що по раю ходив, як повіяв денний холодок. І сховався Адам і його жінка від Господа Бога серед дерев раю.
GEN|3|9|І закликав Господь Бог до Адама, і до нього сказав: Де ти?
GEN|3|10|А той відповів: Почув я Твій голос у раю і злякався, бо нагий я, і сховався.
GEN|3|11|І промовив Господь: Хто сказав тобі, що ти нагий? Чи ти не їв з того дерева, що Я звелів був тобі, щоб ти з нього не їв?
GEN|3|12|А Адам відказав: Жінка, що дав Ти її, щоб зо мною була, вона подала мені з того дерева, і я їв.
GEN|3|13|Тоді Господь Бог промовив до жінки: Що це ти наробила? А жінка сказала: Змій спокусив мене, і я їла.
GEN|3|14|І до змія сказав Господь Бог: За те, що зробив ти оце, то ти проклятіший над усю худобу, і над усю звірину польову! На своїм череві будеш плазувати, і порох ти їстимеш у всі дні свойого життя.
GEN|3|15|І Я покладу ворожнечу між тобою й між жінкою, між насінням твоїм і насінням її. Воно зітре тобі голову, а ти будеш жалити його в п'яту.
GEN|3|16|До жінки промовив: Помножуючи, помножу терпіння твої та болі вагітности твоєї. Ти в муках родитимеш діти, і до мужа твого пожадання твоє, а він буде панувати над тобою.
GEN|3|17|І до Адама сказав Він: За те, що ти послухав голосу жінки своєї та їв з того дерева, що Я наказав був тобі, говорячи: Від нього не їж, проклята через тебе земля! Ти в скорботі будеш їсти від неї всі дні свойого життя.
GEN|3|18|Тернину й осот вона буде родити тобі, і ти будеш їсти траву польову.
GEN|3|19|У поті свойого лиця ти їстимеш хліб, аж поки не вернешся в землю, бо з неї ти взятий. Бо ти порох, і до пороху вернешся.
GEN|3|20|І назвав Адам ім'я своїй жінці: Єва, бо вона була мати всього живого.
GEN|3|21|І зробив Господь Бог Адамові та жінці його одежу шкуряну і зодягнув їх.
GEN|3|22|І сказав Господь Бог: Ось став чоловік, немов один із Нас, щоб знати добро й зло. А тепер коли б не простяг він своєї руки, і не взяв з дерева життя, і щоб він не з'їв, і не жив повік віку.
GEN|3|23|І вислав його Господь Бог із еденського раю, щоб порати землю, з якої узятий він був.
GEN|3|24|І вигнав Господь Бог Адама. А на схід від еденського раю поставив Херувима і меча полум'яного, який обертався навколо, щоб стерегти дорогу до дерева життя.
GEN|4|1|І пізнав Адам Єву, жінку свою, і вона завагітніла, і породила Каїна, і сказала: Набула чоловіка від Господа.
GEN|4|2|А далі вона породила брата йому Авеля. І був Авель пастух отари, а Каїн був рільник.
GEN|4|3|І сталось по деякім часі, і приніс Каїн Богові жертву від плоду землі.
GEN|4|4|А Авель, він також приніс від своїх перворідних з отари та від їхнього лою. І зглянувся Господь на Авеля й на жертву його,
GEN|4|5|а на Каїна й на жертву його не зглянувся. І сильно розгнівався Каїн, і обличчя його похилилось.
GEN|4|6|І сказав Господь Каїнові: Чого ти розгнівався, і чого похилилось обличчя твоє?
GEN|4|7|Отож, коли ти добре робитимеш, то підіймеш обличчя своє, а коли недобре, то в дверях гріх підстерігає. І до тебе його пожадання, а ти мусиш над ним панувати.
GEN|4|8|І говорив Каїн до Авеля, брата свого. І сталось, як були вони в полі, повстав Каїн на Авеля, брата свого, і вбив його.
GEN|4|9|І сказав Господь Каїнові: Де Авель, твій брат? А той відказав: Не знаю. Чи я сторож брата свого?
GEN|4|10|І сказав Господь: Що ти зробив? Голос крови брата твого взиває до Мене з землі.
GEN|4|11|А тепер ти проклятий від землі, що розкрила уста свої, щоб прийняти кров твого брата з твоєї руки.
GEN|4|12|Коли будеш ти порати землю, вона більше не дасть тобі сили своєї. Мандрівником та заволокою будеш ти на землі.
GEN|4|13|І сказав Каїн до Господа: Більший мій гріх, аніж можна знести.
GEN|4|14|Ось Ти виганяєш сьогодні мене з цієї землі, і я буду ховатись від лиця Твого. І я стану мандрівником та заволокою на землі, і буде, кожен, хто стріне мене, той уб'є мене.
GEN|4|15|І промовив до нього Господь: Через те кожен, хто вб'є Каїна, семикратно буде пімщений. І вмістив Господь знака на Каїні, щоб не вбив його кожен, хто стріне його.
GEN|4|16|І вийшов Каїн з-перед лиця Господнього, й осів у країні Нод, на схід від Едену.
GEN|4|17|І Каїн пізнав свою жінку, і стала вона вагітна, і вродила Еноха. І збудував він місто, і назвав ім'я тому містові, як ім'я свого сина: Енох.
GEN|4|18|І народився в Еноха Ірад, а Ірад породив Мехуяїла, а Мехуяїл породив Метушаїла, а Метушаїл породив Ламеха.
GEN|4|19|І взяв собі Ламех дві жінки, ім'я одній Ада, а ймення другій Цілла.
GEN|4|20|І породила Ада Явала, він був батьком тих, що сидять по наметах і мають череду.
GEN|4|21|А ймення брата його Ювал, він був батьком усім, хто держить у руках гусла й сопілку.
GEN|4|22|А Цілла також породила Тувалкаїна, що кував всіляку мідь та залізо. А сестра Тувалкаїнова Ноема.
GEN|4|23|І промовив Ламех до жінок своїх: Адо й Цілло, послухайте ви мого голосу, жони Ламехові, почуйте ви слова мого! Бо якби я мужа забив за уразу свою, а дитину за рану свою,
GEN|4|24|і як буде усемеро пімщений Каїн, то Ламех у сімдесятеро й семеро!
GEN|4|25|І пізнав Адам ще свою жінку, і сина вона породила. І назвала ймення йому: Сиф, бо Бог дав мені інше насіння за Авеля, що забив його Каїн.
GEN|4|26|А Сифові теж народився був син, і він назвав імення йому: Енош. Тоді зачали були призивати Ймення Господнє.
GEN|5|1|Оце книга нащадків Адамових. Того дня, як створив Бог людину, Він її вчинив на подобу Божу.
GEN|5|2|Чоловіком і жінкою Він їх створив, і поблагословив їх. І того дня, як були вони створені, назвав Він їхнє ймення: Людина.
GEN|5|3|І жив Адам сто літ і тридцять, та й сина породив за подобою своєю та за образом своїм, і назвав ім'я йому: Сиф.
GEN|5|4|І було Адамових днів по тому, як він Сифа породив, вісім сотень літ. І породив він синів і дочок.
GEN|5|5|А всіх Адамових днів було, які жив, дев'ять сотень літ і тридцять літ. Та й помер він.
GEN|5|6|І жив Сиф сто літ і п'ять літ, та й породив він Еноша.
GEN|5|7|І жив Сиф по тому, як Еноша породив, вісім сотень літ і сім літ. І породив він синів і дочок.
GEN|5|8|А були всі дні Сифові дев'ять сотень літ і дванадцять літ.
GEN|5|9|І жив Енош дев'ятдесят літ, та й породив він Кенана.
GEN|5|10|І жив Енош по тому, як Кенана породив, вісім сотень літ і п'ятнадцять літ. І породив він синів та дочок.
GEN|5|11|А були всі Еношеві дні дев'ять сотень літ і п'ять літ. Та й помер він.
GEN|5|12|І жив Кенан сімдесят літ, та й породив він Магалал'їла.
GEN|5|13|І жив Кенан по тому, як породив Магалал'їла, вісім сотень літ і сорок літ. І породив він синів та дочок.
GEN|5|14|А всіх Кенанових днів було дев'ять сотень літ і дев'ять літ. Та й помер він.
GEN|5|15|І жив Магалал'їл шістдесят літ і п'ять літ, та й породив він Яреда.
GEN|5|16|І жив Магалал'їл по тому, як Яреда породив, вісім сотень літ і тридцять літ. І породив він синів та дочок.
GEN|5|17|А були всі дні Магалал'їлові вісім сотень літ і дев'ятдесят і п'ять літ. Та й помер він.
GEN|5|18|І жив Яред сто літ і шістдесят і два роки, та й породив він Еноха.
GEN|5|19|І жив Яред по тому, як породив він Еноха, вісім сотень літ. І породив він синів та дочок.
GEN|5|20|А були всі Яредові дні дев'ять сотень літ і шістдесят і два роки. Та й помер він.
GEN|5|21|І жив Енох шістдесят і п'ять літ, та й породив Метушалаха.
GEN|5|22|І ходив Енох з Богом по тому, як породив він Метушалаха, три сотні літ. І породив він синів та дочок.
GEN|5|23|А всіх Енохових днів було три сотні літ і шістдесят і п'ять літ.
GEN|5|24|І ходив із Богом Енох, і не стало його, бо забрав його Бог.
GEN|5|25|І жив Метушалах сто літ і сімдесят і сім літ, та й Ламеха породив.
GEN|5|26|І жив Метушалах по тому, як породив він Ламеха, сім сотень літ і вісімдесят і два роки. І породив він синів та дочок.
GEN|5|27|А всіх Метушалахових днів було дев'ять сотень літ і шістдесят і дев'ять літ. Та й помер він.
GEN|5|28|І жив Ламех сто літ і вісімдесят і два роки, та й сина породив,
GEN|5|29|ім'я йому назвав: Ной, говорячи: Цей нас потішить у наших ділах та в труді рук наших коло землі, що Господь її викляв.
GEN|5|30|І жив Ламех по тому, як Ноя породив, п'ять сотень літ і дев'ятдесят і п'ять літ. І породив він синів та дочок.
GEN|5|31|А всіх Ламехових днів було сім сотень літ і сімдесят і сім літ. Та й помер він.
GEN|5|32|І був Ной віку п'ять сотень літ, та й породив Ной Сима, Хама та Яфета.
GEN|6|1|І сталося, що розпочала людина розмножуватись на поверхні землі, і їм народилися дочки.
GEN|6|2|І побачили Божі сини людських дочок, що вродливі вони, і взяли собі жінок із усіх, яких вибрали.
GEN|6|3|І промовив Господь: Не буде Мій Дух перемагатися в людині навіки, бо блудить вона. Вона тіло, і дні її будуть сто і двадцять літ.
GEN|6|4|За тих днів на землі були велетні, а також по тому, як стали приходити Божі сини до людських дочок. І вони їм народжували, то були силачі, що славні від віку.
GEN|6|5|І бачив Господь, що велике розбещення людини на землі, і ввесь нахил думки серця її тільки зло повсякденно.
GEN|6|6|І пожалкував був Господь, що людину створив на землі. І засмутився Він у серці Своїм.
GEN|6|7|І промовив Господь: Зітру Я людину, яку Я створив, з поверхні землі, від людини аж до скотини, аж до плазунів, і аж до птаства небесного. Бо жалкую, що їх Я вчинив.
GEN|6|8|Але Ной знайшов милість у Господніх очах.
GEN|6|9|Це ось оповість про Ноя. Ной був чоловік праведний і невинний у своїх поколіннях. Ной з Богом ходив.
GEN|6|10|І Ной породив трьох синів: Сима, Хама й Яфета.
GEN|6|11|І зіпсулась земля перед Божим лицем, і наповнилась земля насильством.
GEN|6|12|І бачив Бог землю, і ось зіпсулась вона, кожне бо тіло зіпсуло дорогу свою на землі.
GEN|6|13|І промовив Господь до Ноя: Прийшов кінець кожному тілу перед лицем Моїм, бо наповнилась земля насильством від них. І ось Я винищу їх із землі.
GEN|6|14|Зроби собі ковчега з дерева ґофер. З перегородками зробиш ковчега, і смолою осмолиш його ізсередини та ізнадвору.
GEN|6|15|І отак його зробиш: три сотні ліктів довжина ковчега, п'ятдесят ліктів ширина йому, а тридцять ліктів височина йому.
GEN|6|16|Отвір учиниш в ковчезі, і звузиш на лікоть його від гори, а вхід до ковчегу влаштуєш на боці його. Зробиш його на поверхи долішні, другорядні й третьорядні.
GEN|6|17|А Я ось наведу потоп, воду на землю, щоб з-під неба винищити кожне тіло, що в ньому дух життя. Помре все, що на землі!
GEN|6|18|І складу Я заповіта Свойого з тобою, і ввійдеш до ковчегу ти, і сини твої, і жінка твоя, і жінки твоїх синів із тобою.
GEN|6|19|І впровадиш до ковчегу по двоє з усього, з усього живого, із кожного тіла, щоб їх заховати живими з тобою. Вони будуть самець і самиця.
GEN|6|20|Із птаства за родом його, і з худоби за родом її, і з усіх плазунів на землі за родом їх, по двоє з усього увійдуть до тебе, щоб їх зберегти живими.
GEN|6|21|А ти набери собі з кожної їжі, що вона на споживання, і буде для тебе й для них на поживу.
GEN|6|22|І зробив Ной усе, як звелів йому Бог, так зробив він.
GEN|7|1|І сказав Господь Ноєві: Увійди ти й увесь дім твій до ковчегу, бо Я бачив тебе праведним перед лицем Своїм в оцім роді.
GEN|7|2|Із усякої чистої худоби візьмеш собі по семеро, самця та самицю її, а з худоби нечистої двоє: самця та самицю її.
GEN|7|3|Також із птаства небесного по семеро, самця та самицю, щоб насіння сховати живим на поверхні всієї землі.
GEN|7|4|Ось бо по семи днях Я литиму на землю дощ сорок день і сорок ночей, і всяку істоту, яку Я вчинив, зітру з-над поверхні землі!
GEN|7|5|І зробив Ной усе, як звелів був Господь.
GEN|7|6|А Ной був віку шостисот літ, і стався потоп, вода на землі.
GEN|7|7|І ввійшов Ной, і сини його, і жінка його, і невістки його з ним до ковчегу перед водою потопу.
GEN|7|8|Із чистої худоби та з худоби, що нечиста вона, і з птаства, і всього, що плазує на землі,
GEN|7|9|по двоє ввійшли до Ноя до ковчегу, самець і самиця, як Бог Ноєві був ізвелів.
GEN|7|10|І сталося по семи днях, і води потопу линули на землю.
GEN|7|11|Року шостої сотні літ життя Ноєвого, місяця другого, сімнадцятого дня місяця, цього дня відкрилися всі джерела великої безодні, і розчинилися небесні розтвори.
GEN|7|12|І був дощ на землі сорок день і сорок ночей.
GEN|7|13|Того саме дня до ковчегу ввійшов Ной, і Сим, і Хам та Яфет, сини Ноєві, і жінка Ноєва, і три невістки його з ними,
GEN|7|14|вони та всяка звірина за родом її, і всяка худоба за родом її, і всяке плазуюче, що плазує по землі, за родом його, і всяке птаство за родом його, усяка пташка крилата.
GEN|7|15|І ввійшли до Ноя, до ковчегу по двоє із кожного тіла, що в нім дух життя.
GEN|7|16|А те, що ввійшло, самець і самиця з кожного тіла ввійшли, як звелів йому Бог. І замкнув Господь за ним ковчега.
GEN|7|17|І був потоп сорок день на землі, і збільшилась вода, і понесла ковчега. І він високо став над землею.
GEN|7|18|І прибула вода, і сильно збільшилась вона на землі, і пливав ковчег на поверхні води.
GEN|7|19|І дуже-дуже вода на землі прибула, і покрились усі гори високі, що під небом усім.
GEN|7|20|На п'ятнадцять ліктів угору вода прибула, і покрилися гори.
GEN|7|21|І вимерло всяке тіло, що рухається на землі: серед птаства, і серед скотини, і серед звірини, і серед усіх плазунів, що плазують по землі, і кожна людина.
GEN|7|22|Усе, що в ніздрях його дух життя, з усього, що на суходолі вимерло було.
GEN|7|23|І винищив Бог усяку істоту на поверхні землі, від людини аж до скотини, аж до плазуна, і аж до птаства небесного, вони стерлись з землі. І зостався тільки Ной та те, що з ним у ковчезі було.
GEN|7|24|І прибувала вода на землі сто і п'ятдесят день.
GEN|8|1|І згадав Бог про Ноя, і про кожну звірину та про всяку худобу, що були з ним у ковчезі. І Бог навів вітра на землю, і вода заспокоїлась.
GEN|8|2|І закрились джерела безодні та небесні розтвори, і дощ з неба спинився.
GEN|8|3|І верталась вода з-над землі, верталась постійно. І стала вода спадати по ста й п'ятидесяти днях.
GEN|8|4|А сьомого місяця, на сімнадцятий день місяця ковчег спинився на горах Араратських.
GEN|8|5|І постійно вода спадала аж до десятого місяця. А першого дня десятого місяця завиднілися гірські вершки.
GEN|8|6|І сталося по сорока днях, Ной відчинив вікно ковчегу, що його він зробив.
GEN|8|7|І вислав він крука. І літав той туди та назад, аж поки не висохла вода з-над землі.
GEN|8|8|І послав він від себе голубку, щоб побачити, чи не спала вода з-над землі.
GEN|8|9|Та не знайшла та голубка місця спочинку для стопи своєї ноги, і вернулась до нього до ковчегу, бо стояла вода на поверхні всієї землі. І вистромив руку, і взяв він її, та й до себе в ковчег упустив її.
GEN|8|10|І він зачекав іще других сім день, і знову з ковчегу голубку послав.
GEN|8|11|І голубка вернулась до нього вечірнього часу, і ось у неї в дзюбку лист оливковий зірваний. І довідався Ной, що спала вода з-над землі.
GEN|8|12|І він зачекав іще других сім день, і голубку послав. І вже більше до нього вона не вернулась.
GEN|8|13|І сталося, року шістсотого й першого, місяця першого, першого дня місяця висохла вода з-над землі. І Ной зняв даха ковчегу й побачив: аж ось висохла поверхня землі!
GEN|8|14|А місяця другого, двадцятого й сьомого дня місяця висохла земля.
GEN|8|15|І промовив Ноєві Господь, кажучи:
GEN|8|16|Вийди з ковчегу ти, а з тобою жінка твоя, і сини твої, і невістки твої.
GEN|8|17|Кожну звірину, що з тобою вона, від кожного тіла з-посеред птаства, і з-посеред скотини, і з-посеред усіх плазунів, що плазують по землі, повиводь із собою. І хай рояться вони на землі, і нехай на землі вони плодяться та розмножуються.
GEN|8|18|І вийшов Ной, а з ним сини його, і жінка його, і невістки його.
GEN|8|19|Кожна звірина, кожен плазун, усе птаство, усе, що рухається на землі, за родами їхніми вийшли з ковчегу вони.
GEN|8|20|І збудував Ной жертівника Господеві. І взяв він із кожної чистої худоби й з кожного чистого птаства, і приніс на жертівнику цілопалення.
GEN|8|21|І почув Господь пахощі любі, і в серці Своєму промовив: Я вже більше не буду землі проклинати за людину, бо нахил людського серця лихий від віку його молодого. І вже більше не вбиватиму всього живого, як то Я вчинив був.
GEN|8|22|Надалі, по всі дні землі, сівба та жнива, і холоднеча та спека, і літо й зима, і день та ніч не припиняться!
GEN|9|1|І поблагословив Бог Ноя й синів його, та й промовив: Плодіться й розмножуйтеся, та наповнюйте землю!
GEN|9|2|І ляк перед вами, і страх перед вами буде між усією звіриною землі, і між усім птаством небесним, між усім, чим роїться земля, і між усіма рибами моря. У ваші руки віддані вони.
GEN|9|3|Усе, що плазує, що живе воно, буде вам на їжу. Як зелену ярину Я віддав вам усе.
GEN|9|4|Тільки м'яса з душею його, цебто з кров'ю його, не будете ви споживати.
GEN|9|5|А тільки Я буду жадати вашу кров із душ ваших, з руки кожної звірини буду жадати її, і з руки чоловіка, з руки кожного брата його Я буду жадати душу людську.
GEN|9|6|Хто виллє кров людську з людини, то виллята буде його кров, бо Він учинив людину за образом Божим.
GEN|9|7|Ви ж плодіться й розмножуйтеся, роїться на землі та розмножуйтесь на ній!
GEN|9|8|І сказав Бог до Ноя та до синів його з ним, кажучи:
GEN|9|9|А Я, ось Свого заповіта укладаю Я з вами та з вашим потомством по вас.
GEN|9|10|І з кожною живою душею, що з вами: серед птаства, серед худоби, і серед усієї земної звірини з вами, від усіх, що виходять з ковчегу, до всієї земної звірини.
GEN|9|11|І Я укладу заповіта Свого з вами, і жодне тіло не буде вже знищене водою потопу, і більш не буде потопу, щоб землю нищити.
GEN|9|12|І Бог промовляв: Оце знак заповіту, що даю Я його поміж Мною та вами, і поміж кожною живою душею, що з вами, на вічні покоління:
GEN|9|13|Я веселку Свою дав у хмарі, і стане вона за знака заповіту між Мною та між землею.
GEN|9|14|І станеться, коли над землею Я хмару захмарю, то буде виднітися в хмарі веселка.
GEN|9|15|І згадаю про Свого заповіта, що між Мною й між вами, і між кожною живою душею в кожному тілі. І більш не буде вода для потопу, щоб вигубляти кожне тіло.
GEN|9|16|І буде веселка у хмарі, і побачу її, щоб пам'ятати про вічний заповіт між Богом і між кожною живою душею в кожному тілі, що воно на землі.
GEN|9|17|І сказав Бог до Ноя: Це знак заповіту, що Я встановив поміж Мною й поміж кожним тілом, що воно на землі.
GEN|9|18|І були сини Ноєві, що вийшли з ковчегу: Сим, і Хам, і Яфет. А Хам він був батько Ханаанів.
GEN|9|19|Оці троє були сини Ноєві, і від них залюднилася вся земля.
GEN|9|20|І зачав був Ной, муж землі, садити виноград.
GEN|9|21|І пив він вино та й упився, й обнажився в середині свого намету.
GEN|9|22|І побачив Хам, батько Ханаанів, наготу батька свого, та й розказав обом браттям своїм надворі.
GEN|9|23|Узяли тоді Сим та Яфет одежину, і поклали обидва на плечі свої, і позадкували, та й прикрили наготу батька свого. Вони відвернули дозаду обличчя свої, і не бачили наготи батька свого.
GEN|9|24|А Ной витверезився від свого вина, і довідався, що йому був учинив його син наймолодший.
GEN|9|25|І сказав він: Проклятий будь Ханаан, він буде рабом рабів своїм браттям!
GEN|9|26|І сказав він: Благословенний Господь, Симів Бог, і хай Ханаан рабом буде йому!
GEN|9|27|Нехай Бог розпросторить Яфета, і нехай пробуває в наметах він Симових, і нехай Ханаан рабом буде йому!
GEN|9|28|А Ной жив по потопі триста літ і п'ятдесят літ.
GEN|9|29|А всіх Ноєвих днів було дев'ятсот літ і п'ятдесят літ. Та й помер.
GEN|10|1|Оце нащадки синів Ноєвих: Сима, Хама та Яфета. А їм народились сини по потопі:
GEN|10|2|Сини Яфетові: Ґомер, і Маґоґ, і Мадай, і Яван, і Тувал, і Мешех, і Тирас.
GEN|10|3|А сини Ґомерові: Ашкеназ, і Рифат, і Тоґарма.
GEN|10|4|А сини Явана: Еліша, і Таршіш, і китти, і додани.
GEN|10|5|Від них відділилися острови народів у їхніх краях, кожний за мовою своєю, за своїми родами, у народах своїх.
GEN|10|6|А сини Хамові: Куш, і Міцраїм, і Фут, і Ханаан.
GEN|10|7|А сини Кушові: Сева, і Хавіла, і Савта, і Раама, і Савтеха. А сини Раами: Шева та Дедан.
GEN|10|8|Куш же породив Німрода, він розпочав на землі велетнів.
GEN|10|9|Він був дужий мисливець перед Господнім лицем. Тому то говориться: Як Німрод, дужий мисливець перед Господнім лицем.
GEN|10|10|А початком царства його були: Вавилон, і Ерех, і Аккад, і Калне в землі Шінеар.
GEN|10|11|З того краю вийшов Ашшур, та й збудував Ніневію, і Реховот-Ір, і Калах,
GEN|10|12|і Ресен поміж Ніневією та поміж Калахом, він оте місто велике.
GEN|10|13|А Міцраїм породив лудів, і анамів, і легавів, і нафтухів,
GEN|10|14|і патрусів, і каслухів, що звідси пішли филистимляни, і кафторів.
GEN|10|15|А Ханаан породив Сидона, свого перворідного, та Хета,
GEN|10|16|і Евусеянина, і Амореянина, і Ґірґашеянина,
GEN|10|17|і Хіввеянина, і Аркеянина, і Синеянина,
GEN|10|18|і Арвадеянина, і Цемареянина, і Хаматеянина. А потім розпорошилися роди Ханаанеянина.
GEN|10|19|І була границя Ханаанеянина від Сидону в напрямі аж до Ґерару, аж до Ґази, у напрямі аж до Содому, і до Гомори, і до Адми, і до Цевоїму, аж до Лашу.
GEN|10|20|Оце сини Хамові, за їхніми родами, за мовами їхніми, у їхніх країнах, у їхніх народах.
GEN|10|21|А Симові теж народились йому, він батько всіх синів Еверових, брат старший Яфетів.
GEN|10|22|Сини Симові: Елам, і Ашшур, і Арпахшад, і Луд, і Арам.
GEN|10|23|А Арамові сини: Уц, і Хул, і Ґетер, і Маш.
GEN|10|24|А Арпахшад породив Шелаха, а Шелах породив Евера.
GEN|10|25|А Еверові народилося двоє синів: ім'я першому Пелеґ, бо за днів його поділилась земля, а ймення його брата Йоктан.
GEN|10|26|А Йоктан породив Алмодада, і Шелефа, і Хасар-Мавета, і Єраха,
GEN|10|27|і Гадорама, і Узала, і Диклу,
GEN|10|28|і Увала, і Авімаїла, і Шеву,
GEN|10|29|і Офіра, і Хавілу, і Йовава. Усі вони сини Йоктанові.
GEN|10|30|А оселя їхня була від Меші в напрямі аж до Сефару, гори східньої.
GEN|10|31|Оце сини Симові, за їхніми родами, за мовами їхніми, у їхніх країнах, у їхніх народах.
GEN|10|32|Оце роди синів Ноєвих, за нащадками їхніми, у їхніх народах. І народи від них поділились на землі по потопі.
GEN|11|1|І була вся земля одна мова та слова одні.
GEN|11|2|І сталось, як рушали зо Сходу вони, то в Шинеарському краї рівнину знайшли, і оселилися там.
GEN|11|3|І сказали вони один одному: Ану, наробімо цегли, і добре її випалімо! І сталася цегла для них замість каменя, а смола земляна була їм за вапно.
GEN|11|4|І сказали вони: Тож місто збудуймо собі, та башту, а вершина її аж до неба. І вчинімо для себе ймення, щоб ми не розпорошилися по поверхні всієї землі.
GEN|11|5|І зійшов Господь, щоб побачити місто та башту, що людські сини будували її.
GEN|11|6|І промовив Господь: Один це народ, і мова одна для всіх них, а це ось початок їх праці. Не буде тепер нічого для них неможливого, що вони замишляли чинити.
GEN|11|7|Тож зійдімо, і змішаймо там їхні мови, щоб не розуміли вони мови один одного.
GEN|11|8|І розпорошив їх звідти Господь по поверхні всієї землі, і вони перестали будувати те місто.
GEN|11|9|І тому то названо ймення йому: Вавилон, бо там помішав Господь мову всієї землі. І розпорошив їх звідти Господь по поверхні всієї землі.
GEN|11|10|Оце нащадки Симові: Сим був віку ста літ, та й породив Арпахшада, два роки по потопі.
GEN|11|11|І жив Сим по тому, як породив Арпахшада, п'ять сотень літ. І породив він синів і дочок.
GEN|11|12|А Арпахшад жив тридцять і п'ять літ, та й породив він Шелаха.
GEN|11|13|І жив Арпахшад по тому, як породив він Шелаха, чотири сотні літ та три роки. І породив він синів та дочок.
GEN|11|14|Шелах же жив тридцять літ, та й породив він Евера.
GEN|11|15|І жив Шелах по тому, як породив він Евера, чотири сотні літ і три роки. І породив він синів та дочок.
GEN|11|16|Евер же жив тридцять літ і чотири, та й породив він Пелеґа.
GEN|11|17|І жив Евер по тому, як породив він Пелеґа, чотири сотні літ і тридцять літ. І породив він синів та дочок.
GEN|11|18|Пелеґ же жив тридцять літ, та й породив Реу.
GEN|11|19|І жив Пелеґ по тому, як породив Реу, дві сотні літ і дев'ять літ. І породив він синів та дочок.
GEN|11|20|А Реу жив тридцять і два роки, та й породив Серуґа.
GEN|11|21|І жив Реу по тому, як породив Серуґа, дві сотні літ і сім літ. І породив він синів та дочок.
GEN|11|22|А Серуґ жив тридцять літ, та й породив Нахора.
GEN|11|23|І жив Серуґ по тому, як породив Нахора, дві сотні літ. І породив він синів та дочок.
GEN|11|24|А Нахор жив двадцять літ і дев'ять, та й породив він Тераха.
GEN|11|25|І жив Нахор по тому, як породив він Тераха, сотню літ і дев'ятнадцять літ. І породив він синів та дочок.
GEN|11|26|Терах же жив сімдесят літ, та й породив Аврама, і Нахора, і Гарана.
GEN|11|27|А оце нащадки Терахові: Терах породив Аврама, і Нахора, і Гарана. А Гаран породив Лота.
GEN|11|28|Гаран же помер за життя свого батька, у краї свого народження, в Урі халдейському.
GEN|11|29|І побрали Аврам та Нахор для себе жінок. Ім'я Аврамовій жінці Сара, а ймення Нахоровій жінці Мілка, дочка Гарана, Мілчиного батька і батька Їски.
GEN|11|30|А Сара неплідна була, не мала нащадка вона.
GEN|11|31|І взяв Терах Аврама, сина свого, і Лота, сина Гаранового, сина свого сина, і Сару, невістку свою, жінку Аврама, свого сина, та й вийшов з ними з Уру халдейського, щоб піти до краю ханаанського. І прийшли вони аж до Харану, та й там оселилися.
GEN|11|32|І було днів Терахових дві сотні літ та п'ять літ. І Терах помер у Харані.
GEN|12|1|І промовив Господь до Аврама: Вийди зо своєї землі, і від родини своєї, і з дому батька свого до Краю, який Я тобі покажу.
GEN|12|2|І народом великим тебе Я вчиню, і поблагословлю Я тебе, і звеличу ймення твоє, і будеш ти благословенням.
GEN|12|3|І поблагословлю, хто тебе благословить, хто ж тебе проклинає, того прокляну. І благословляться в тобі всі племена землі!
GEN|12|4|І відправивсь Аврам, як сказав був до нього Господь, і з ним пішов Лот. Аврам же мав віку сімдесят літ і п'ять літ, як виходив з Харану.
GEN|12|5|І Аврам узяв Сару, свою жінку, та Лота, сина брата свого, і ввесь маєток, який набули, і людей, що їх набули у Харані, та й вийшли, щоб піти до Краю ханаанського. І до Краю ханаанського вони прибули.
GEN|12|6|І пройшов Аврам по Краю аж до місця Сихему, аж до дуба Мамре. А ханаанеянин тоді проживав у цім Краї.
GEN|12|7|І Господь явився Авраму й сказав: Я дам оцей Край потомству твоєму. І він збудував там жертівника Господеві, що явився йому.
GEN|12|8|А звідти він рушив на гору від сходу від Бет-Елу, і намета свого розіп'яв, Бет-Ел від заходу, а Гай від сходу. І він збудував там Господу жертівника, і прикликав Господнє Ймення.
GEN|12|9|І подавався Аврам усе далі на південь.
GEN|12|10|І стався був голод у Краї. І зійшов Аврам до Єгипту, щоб там перебути, бо голод у Краї тяжкий став.
GEN|12|11|І сталося, як він близько прийшов до Єгипту, то сказав був до жінки своєї Сари: Отож то я знаю, що ти жінка вродлива з обличчя.
GEN|12|12|І станеться, як побачать тебе єгиптяни й скажуть: Це жінка його, то вони мене вб'ють, а тебе позоставлять живою.
GEN|12|13|Скажи ж, що сестра моя ти, щоб добре було через тебе мені, і щоб я позостався живий через тебе.
GEN|12|14|І сталось, як прийшов був Аврам до Єгипту, то єгиптяни побачили жінку, що дуже вродлива вона.
GEN|12|15|І побачили її вельможі фараонові, і хвалили її перед фараоном. І взята була та жінка до дому фараонового.
GEN|12|16|І він для Аврама добро вчинив через неї. І одержав він дрібну та велику худобу, і осли, і раби, і невільниці, і ослиці, верблюди.
GEN|12|17|І вдарив Господь фараона та дім його великими поразами через Сару, Аврамову жінку.
GEN|12|18|І прикликав фараон Аврама й сказав: Що ж то мені ти вчинив? Чому не сказав мені, що вона твоя жінка?
GEN|12|19|Для чого сказав ти: Вона моя сестра? І я собі взяв був за жінку її. А тепер ось жінка твоя, візьми та й іди!
GEN|12|20|І фараон наказав людям про нього. І вислали його, і жінку його, і все, що в нього було.
GEN|13|1|І піднявся Аврам із Єгипту, сам, і жінка його, і все, що в нього було, і Лот разом із ним, до Неґеву.
GEN|13|2|А Аврам був вельми багатий на худобу, на срібло й на золото.
GEN|13|3|І пішов він в мандрівки свої від Неґеву аж до Бет-Елу, аж до місця, де напочатку намет його був поміж Бет-Елом і поміж Гаєм,
GEN|13|4|до місця жертівника, що його він зробив там напочатку. І Аврам там прикликав Господнє Ймення.
GEN|13|5|Так само й у Лота, що з Аврамом ходив, дрібна та велика худоба була та намети.
GEN|13|6|І не вміщала їх та земля, щоб їм разом пробувати, бо великий був їхній маєток, і не могли вони разом пробувати.
GEN|13|7|І сталася сварка поміж пастухами худоби Аврамової та поміж пастухами худоби Лотової. А ханаанеянин та періззеянин сиділи тоді в Краю.
GEN|13|8|І промовив до Лота Аврам: Нехай сварки не буде між мною та між тобою, і поміж пастухами моїми та поміж пастухами твоїми, бо близька ми рідня.
GEN|13|9|Хіба не ввесь Край перед обличчям твоїм? Відділися від мене! Коли підеш ліворуч, то я піду праворуч, а як ти праворуч, то піду я ліворуч.
GEN|13|10|І звів Лот свої очі, і побачив усю околицю Йорданську, що наводнена вся вона аж до Цоару, перед тим, як Содом та Гомору був знищив Господь, як Господній, садок, як єгипетський край!
GEN|13|11|І Лот вибрав собі всю околицю йорданську. І Лот рушив на схід, і вони розлучилися один від одного.
GEN|13|12|Аврам оселився в землі ханаанській, а Лот оселився в рівнинних містах околиці, і наметував аж до Содому.
GEN|13|13|А люди содомські були дуже злі та грішні перед Господом.
GEN|13|14|І промовив Господь до Аврама, коли Лот розлучився із ним: Зведи очі свої, та поглянь із місця, де ти, на північ, і на південь, і на схід, і на захід,
GEN|13|15|бо всю цю землю, яку бачиш, Я її дам навіки тобі та потомству твоєму.
GEN|13|16|І вчиню Я потомство твоє, як той порох землі, так, що коли хто потрапить злічити порох земний, то теж і потомство твоє перелічене буде.
GEN|13|17|Устань, пройдись по Краю вздовж його та вширшки його, бо тобі його дам!
GEN|13|18|І Аврам став наметувати, і прибув, і осів між дубами Мамре, що в Хевроні вони. І він збудував там жертівника Господеві.
GEN|14|1|І сталось за днів Амрафела, царя Шинеару, Арйоха, царя Елласару, Кедор-Лаомера, царя Еламу, і Тидала, царя Ґоїму,
GEN|14|2|вони вчинили війну з Бераєм, царем Содому, і з Біршаєм, царем Гомори, з Шин'авом, царем Адми, і Шемевером, царем Цевоїму, і з царем Белаю, що Цоар тепер.
GEN|14|3|Усі ці зібрались були до долини Сіддім, вона тепер море Солоне.
GEN|14|4|Дванадцять літ служили вони Кедор-Лаомерові, а року тринадцятого повстали.
GEN|14|5|А року чотирнадцятого прибув Кедор-Лаомер та царі, що були з ним, і побили Рефаїв в Аштерот-Карнаїмі, і Зузів у Гамі, і Емів у Шаве-Кір'ятаїмі,
GEN|14|6|і Хорянина в горах Сеїру аж до Ел-Парану, що він при пустині.
GEN|14|7|І вернулись вони, і прибули до Ен-Мішпату, воно тепер Кадеш, і звоювали всю землю Амалика, а також Аморея, що сидів у Хаццон-Тамарі.
GEN|14|8|І вийшов цар Содому, і цар Гомори, і цар Адми, і цар Цевоїму, і цар Белаю, тепер він Цоар, і вишикувалися з ними на бій у долині Сіддім,
GEN|14|9|із Кедор-Лаомером, царем Еламу, і Тидалом, царем Ґоїму, і Амрафелом, царем Шинеару, і Арйохом, царем Елласару, чотири царі проти п'ятьох.
GEN|14|10|А долина Сіддім була повна смоляних ям; і втекли цар Содому й цар Гомори, та й попадали туди, а позосталі повтікали на гору.
GEN|14|11|І взяли вони ввесь маєток Содому й Гомори, і всю їхню поживу, і пішли.
GEN|14|12|І взяли вони Лота, сина брата Аврамового, бо пробував у Содомі, і добро його та й пішли.
GEN|14|13|І прийшов був недобиток, та й розповів єврею Аврамові, а він жив між дубами амореянина Мамре, брата Ешколового й брата Анерового, Аврамових спільників.
GEN|14|14|І почув Аврам, що небіж його взятий у неволю, та й узброїв своїх вправних слуг, що в домі його народились, три сотні й вісімнадцять, і погнався до Дану.
GEN|14|15|І він поділився на гурти вночі, він та раби його, і розбив їх, і гнався за ними аж до Хови, що ліворуч Дамаску.
GEN|14|16|І вернув він усе добро, а також Лота, небожа свого, і добро його повернув, а також жінок та людей.
GEN|14|17|Тоді цар Содому вийшов назустріч йому, як він повертався, розбивши Кедор-Лаомера та царів, що були з ним, до долини Шаве, вона тепер долина Царська.
GEN|14|18|А Мелхиседек, цар Салиму, виніс хліб та вино. А він був священик Бога Всевишнього.
GEN|14|19|І поблагословив він його та й промовив: Благословенний Аврам від Бога Всевишнього, що створив небо й землю.
GEN|14|20|І благословенний Бог Всевишній, що видав у руки твої ворогів твоїх. І Аврам дав йому десятину зо всього.
GEN|14|21|І сказав цар содомський Аврамові: Дай мені людей, а маєток візьми собі.
GEN|14|22|Аврам же сказав цареві содомському: Я звів свою руку до Господа, Бога Всевишнього, Творця неба й землі,
GEN|14|23|що від нитки аж до ремінця сандалів я не візьму з того всього, що твоє, щоб ти не сказав: Збагатив я Аврама.
GEN|14|24|Я не хочу нічого, даси тільки те, що слуги поїли, та частину людям, що зо мною ходили: Анер, Ешкол і Мамре, частину свою вони візьмуть.
GEN|15|1|По цих-о подіях було слово Господнє Аврамові в видінні таке: Не бійся, Авраме, Я тобі щит, нагорода твоя вельми велика.
GEN|15|2|А Аврам відізвався: Господи, Господи, що даси Ти мені, коли я бездітний ходжу, а керівник мого господарства він Елі-Езер із Дамаску.
GEN|15|3|І сказав Аврам: Отож, Ти не дав нащадка мені, і ото мій керівник спадкоємець мені.
GEN|15|4|І ось слово Господнє до нього таке: Він не буде спадкоємець тобі, але той, хто вийде з твойого нутра, він буде спадкоємець тобі.
GEN|15|5|І Господь його вивів надвір та й сказав: Подивися на небо, та зорі злічи, коли тільки потрапиш ти їх полічити. І до нього прорік: Таким буде потомство твоє!
GEN|15|6|І ввірував Аврам Господеві, а Він залічив йому те в праведність.
GEN|15|7|І промовив до нього: Я Господь, що вивів тебе з Уру халдейського, щоб дати тобі землю оцю, щоб став ти спадкоємець її.
GEN|15|8|І промовив Аврам: Господи, Господи, з чого я довідаюся, що буду спадкоємець її?
GEN|15|9|Він же промовив до нього: Візьми трилітнє теля, і трилітню козу, і трилітнього барана, і горлицю, і пташеня голубине.
GEN|15|10|І взяв він для Нього все те, і розсік його пополовині, і дав кожну частину його відповідно до другої, але птаства не розсік.
GEN|15|11|І зліталося хиже птаство на трупи, та Аврам відганяв його.
GEN|15|12|Коли ж сонце схилялось на захід, то спав сон на Аврама. І ось спадає на нього жах темний, великий.
GEN|15|13|І промовив Господь до Аврама: Добре знай, що потомство твоє буде приходьком в землі не своїй. І будуть служити вони, і будуть їх мучити чотири сотні літ.
GEN|15|14|Але народ, якому служити вони будуть, Я засуджу; та вони потім вийдуть з великим маєтком.
GEN|15|15|А ти до своєї рідні прийдеш у мирі, у старості добрій похований будеш.
GEN|15|16|А покоління четверте повернеться сюди, бо досі не повний ще гріх амореянина.
GEN|15|17|І сталось, коли зайшло сонце й була темрява, то ось появилась мов димуюча піч, та смолоскип огняний перейшов поміж тими кусками жертви.
GEN|15|18|І того дня склав Господь заповіта з Аврамом, говорячи: Потомству твоєму Я дав оцю землю від річки Єгипту аж до річки великої, до річки Ефрата:
GEN|15|19|хенеянина, і кенізеянина, і кадмонеянина,
GEN|15|20|і хіттеянина, і періззеянина, і рефаеянина,
GEN|15|21|і амореянина, і ханаанеянина, і ґірґашеянина, і евусеянина.
GEN|16|1|А Сара, Аврамова жінка, не родила йому. І в неї була єгиптянка невільниця, а ймення їй Аґар.
GEN|16|2|І сказала Сара Аврамові: Ось Господь затримав мене від породу. Прийди ж до моєї невільниці, може від неї одержу я сина. І послухався Аврам голосу Сари.
GEN|16|3|І взяла Сара, Аврамова жінка, єгиптянку Аґар, свою невільницю, по десяти літах перебування Аврамового в землі ханаанській, і дала її Аврамові, чоловікові своєму, за жінку.
GEN|16|4|І він увійшов до Аґари, і вона зачала. Як вона ж побачила, що зачала, то стала легковажити господиню свою.
GEN|16|5|І сказала Сара Аврамові: Моя кривда на тобі! Я дала була свою невільницю до лоня твого, а як вона побачила, що зачала, то стала легковажити мене. Нехай розсудить Господь поміж мною та поміж тобою!
GEN|16|6|І промовив Аврам до Сари: Таж невільниця твоя в руці твоїй! Зроби їй те, що вгодне в очах твоїх. І Сара гнобила її. І втекла Аґар від обличчя її.
GEN|16|7|І знайшов її Ангол Господній біля джерела води на пустині, біля джерела на дорозі до Шур,
GEN|16|8|і сказав: Аґаро, Сарина невільнице, звідки ж то прийшла ти, і куди ти йдеш? Та відказала: Я втікаю від обличчя Сари, пані моєї.
GEN|16|9|А Ангол Господній промовив до неї: Вернися до пані своєї, і терпи під руками її!
GEN|16|10|І Ангол Господній промовив до неї: Сильно розмножу потомство твоє, і через безліч буде воно незліченне.
GEN|16|11|І Ангол Господній до неї сказав: Ось ти зачала, і сина породиш, і назвеш ім'я йому Ізмаїл, бо прислухавсь Господь до твоєї недолі.
GEN|16|12|А він буде як дикий осел між людьми, рука його на всіх, а рука всіх на нього. І буде він жити при всіх своїх браттях.
GEN|16|13|І назвала вона Ймення Господа, що мовив до неї: Ти Бог видіння! Бо сказала вона: Чи й тут я дивилась на Того, Хто бачить мене?
GEN|16|14|Тому джерело було назване Джерело Живого, Хто бачить мене, воно поміж Кадешем та поміж Баредом.
GEN|16|15|І вродила Аґар Аврамові сина, а Аврам назвав ім'я свого сина, що вродила Аґар: Ізмаїл.
GEN|16|16|А Аврам був віку восьмидесяти літ і шести літ, коли Аґар вродила була Аврамові Ізмаїла.
GEN|17|1|І був Аврам віку дев'ятидесяти літ і дев'яти літ, коли явився Господь Аврамові та й промовив до нього: Я Бог Всемогутній! Ходи перед лицем Моїм, і будь непорочний!
GEN|17|2|І дам Я Свого заповіта поміж Мною та поміж тобою, і дуже-дуже розмножу тебе.
GEN|17|3|І впав Аврам на обличчя своє, а Бог до нього промовляв, говорячи:
GEN|17|4|Я, ось Мій заповіт із тобою, і станеш ти батьком багатьох народів.
GEN|17|5|І не буде вже кликатись ім'я твоє: Аврам, але буде ім'я твоє: Авраам, бо вчинив Я тебе батьком багатьох народів.
GEN|17|6|І вчиню Я тебе дуже-дуже плідним, і вчиню, щоб вийшли з тебе народи, і царі з тебе вийдуть.
GEN|17|7|І Я складу заповіта Свого поміж Мною та поміж тобою, і поміж твоїм потомством по тобі на їхні покоління на вічний заповіт, що буду Я Богом для тебе й для нащадків твоїх по тобі.
GEN|17|8|І дам Я тобі та потомству твоєму по тобі землю скитання твого, увесь Край ханаанський, на вічне володіння, і Я буду їм Богом.
GEN|17|9|І сказав Авраамові Бог: А ти заповіта Мого стерегтимеш, ти й потомство твої по тобі в їхніх поколіннях.
GEN|17|10|То Мій заповіт, що його ви виконувать будете, поміж Мною й поміж вами, і поміж потомством твоїм по тобі: нехай кожен чоловічої статі буде обрізаний у вас.
GEN|17|11|І будете ви обрізані на тілі крайньої плоті вашої, і стане це знаком заповіту поміж Мною й поміж вами.
GEN|17|12|А кожен чоловічої статі восьмиденний у вас буде обрізаний у всіх ваших поколіннях, як народжений дому, так і куплений за срібло з-поміж чужоплемінних, що він не з потомства твого.
GEN|17|13|Щодо обрізання, нехай буде обрізаний уроджений дому твого й куплений за срібло твоє, і буде Мій заповіт на вашім тілі заповітом вічним.
GEN|17|14|А необрізаний чоловічої статі, що не буде обрізаний на тілі своєї крайньої плоті, то стята буде душа та з народу свого, він зірвав заповіта Мого!
GEN|17|15|І сказав Авраамові Бог: Сара, жінка твоя, нехай свого ймення не кличе вже: Сара, бо ім'я їй: Сарра.
GEN|17|16|І поблагословлю Я її, і теж з неї дам сина тобі. І поблагословлю Я її, і стануться з неї народи, і царі народів будуть із неї.
GEN|17|17|І впав Авраам на обличчя своє, і засміявся. І подумав він у серці своїм: Чи в столітнього буде народжений, і чи Сарра в віці дев'ятидесяти літ уродить?
GEN|17|18|А до Бога сказав Авраам: Хоча б Ізмаїл жив перед лицем Твоїм!
GEN|17|19|Бог же сказав: Але Сарра, твоя жінка, сина породить тобі, а ти назвеш ім'я йому Ісак. І Свого заповіта з ним Я складу, щоб був вічний заповіт для нащадків його по нім.
GEN|17|20|А щодо Ізмаїла, Я послухав тебе: Ось Я поблагословлю його, і вчиню його плідним, і дуже-дуже розмножу його. Він породить дванадцять князів, і великим народом учиню Я його.
GEN|17|21|А Свого заповіта Я складу з Ісаком, що його Сарра вродить тобі на цей час другого року.
GEN|17|22|І Він перестав говорити з ним. І Бог вознісся від Авраама.
GEN|17|23|І взяв Авраам Ізмаїла, сина свого, і всіх уроджених у домі його, і всіх, хто куплений за срібло його, кожного чоловічої статі з-поміж людей Авраамового дому, і обрізав тіло крайньої плоті їх того самого дня, як Бог говорив з ним.
GEN|17|24|А Авраам був віку дев'ятидесяти й дев'яти літ, як обрізано було тіло крайньої плоті його.
GEN|17|25|А Ізмаїл був віку тринадцяти літ, як обрізано було тіло крайньої плоті його.
GEN|17|26|Того самого дня був обрізаний Авраам та Ізмаїл, син його.
GEN|17|27|І всі мужі дому його, народжені дому й куплені за срібло з-поміж чужоплемінних, були обрізані з ним.
GEN|18|1|І явився до нього Господь між дубами Мамре, а він сидів при вході в намет під час денної спеки.
GEN|18|2|І він ізвів очі свої та й побачив: ось три Мужі стоять біля нього. І побачив, і вибіг із входу намету назустріч Їм, і вклонився до землі,
GEN|18|3|та й промовив: Господи, коли тільки знайшов я милість в очах Твоїх, не проходь повз Свойого раба!
GEN|18|4|Принесуть трохи води, і ноги Свої помийте, і спочиньте під деревом.
GEN|18|5|І хай хліба шматок принесу я, а Ви підкріпіть серце Ваше. Потому підете, бо на те Ви йдете повз свойого раба. І сказали вони: Зроби так, як сказав.
GEN|18|6|І Авраам поспішив до намету до Сарри й сказав: Візьми швидко три міри пшеничної муки, заміси, і зроби коржі.
GEN|18|7|І побіг Авраам до товару, і взяв молоде та добре теля, і дав слузі, а той швидко його приготовив.
GEN|18|8|І взяв масла й молока, та теля приготовлене, та й поклав перед Ними, а сам став біля Них під деревом. І їли Вони.
GEN|18|9|І сказали до нього: Де Сарра, жінка твоя? А він відказав: Ось у наметі.
GEN|18|10|І сказав один з Них: Я напевно вернуся до тебе за рік цього самого часу. І ось буде син у Сарри, жінки твоєї... А Сарра це чула при вході намету, що був за Ним.
GEN|18|11|Авраам же та Сарра старі були, віку похилого. У Сарри перестало бувати звичайне жіноче.
GEN|18|12|І засміялася Сарра в нутрі своїм, говорячи: Коли я зів'яла, то як станеться розкіш мені? Таж пан мій старий!
GEN|18|13|І сказав Господь до Авраама: Чого то сміялася Сарра отак: Чи ж справді вроджу, коли я зостарілась?
GEN|18|14|Чи для Господа є річ занадто трудна? На означений час Я вернуся до тебе за рік цього самого часу, Сарра ж тоді матиме сина.
GEN|18|15|А Сарра відріклася, говорячи: Не сміялася я, бо боялась. Але Він відказав: Ні, таки сміялася ти!
GEN|18|16|І повставали звідти ті Мужі, і поглянули на Содом, а Авраам пішов з Ними, щоб Їх відпровадити.
GEN|18|17|А Господь сказав: Чи Я від Авраама втаю, що Я маю зробити?
GEN|18|18|Бож Авраам справді стане народом великим та дужим, і в ньому поблагословляться всі народи землі!
GEN|18|19|Бо вибрав Я його, щоб він наказав синам своїм і домові своєму по собі. І будуть вони дотримуватися дороги Господньої, щоб чинити справедливість та право, а то для того, щоб Господь здійснив на Авраамові, що сказав був про нього.
GEN|18|20|І промовив Господь: Через те, що крик Содому й Гомори великий, і що гріх їхній став дуже тяжкий,
GEN|18|21|зійду ж Я та й побачу, чи не вчинили вони так, як крик про них, що доходить до Мене, тоді їм загибіль, а як ні то побачу.
GEN|18|22|І повернулися звідти ті Мужі, і пішли до Содому, а Авраам усе ще стояв перед Господнім лицем.
GEN|18|23|І Авраам підійшов та й промовив: Чи погубиш також праведного з нечестивим?
GEN|18|24|Може є п'ятдесят праведних у цьому місті, чи також вигубиш і не пробачиш цій місцевості ради п'ятидесяти тих праведних, що в ньому є?
GEN|18|25|Не можна Тобі чинити так, щоб убити праведного з нечестивим, бо стане праведний як нечестивий, цього ж не можна Тобі! Чи ж Той, Хто всю землю судить, не вчинить правди?
GEN|18|26|І промовив Господь: Коли Я в Содомі, у цьому місті, знайду п'ятдесят праведних, то вибачу цілій місцевості ради них.
GEN|18|27|І відповів Авраам та й промовив: Оце я осмілився був говорити до Господа свого, а я порох та попіл.
GEN|18|28|Може п'ятдесят тих праведних не матиме п'яти, чи Ти знищиш ціле місто через п'ятьох? І промовив Господь: Не знищу, коли там знайду сорок і п'ять!
GEN|18|29|І промовив до Нього він ще, та й сказав: Може сорок там знайдеться? А Господь відказав: Не зроблю й ради сорока!
GEN|18|30|І сказав Авраам: Хай не гніває це мого Господа, і нехай я скажу: Може тридцять там знайдеться? А Господь відказав: Не зроблю, коли й тридцять знайду там!
GEN|18|31|І сказав Авраам: Оце я осмілився був говорити до Господа мого: Може двадцять там знайдеться? А Господь відказав: Не зроблю й ради двадцяти!
GEN|18|32|І сказав Авраам: Хай не гніває це мого Господа, і нехай я скажу тільки разу цього: Може хоч десять там знайдеться? А Господь відказав: Не знищу й ради десятьох!
GEN|18|33|І пішов Господь, як скінчив говорити до Авраама. А Авраам вернувся до свого місця.
GEN|19|1|І прибули обидва Анголи до Содому надвечір, а Лот сидів у брамі содомській. І побачив Лот, і встав їм назустріч, і вклонився обличчям до землі,
GEN|19|2|та й промовив: Ось, панове мої, зайдіть до дому вашого раба, і переночуйте, і помийте ноги свої, а рано встанете й підете на дорогу свою. А вони відказали: Ні, бо будемо ми ночувати на вулиці.
GEN|19|3|А він сильно на них налягав, і вони до нього з дороги зійшли, і ввійшли до дому його. І вчинив він для них прийняття, і напік прісного і їли вони.
GEN|19|4|Ще вони не полягали, а люди того міста, люди Содому від малого аж до старого, увесь народ звідусюди оточили той дім.
GEN|19|5|І вони закричали до Лота, і сказали йому: Де ті мужі, що ночі цієї до тебе прийшли? Виведи їх до нас, щоб нам їх пізнати!
GEN|19|6|І Лот вийшов до входу до них, а двері замкнув за собою,
GEN|19|7|і сказав: Браття мої, не чиніть лихого!
GEN|19|8|Ось у мене дві доньки, що мужа не пізнали. Нехай я їх до вас виведу, а ви їм робіть, що вам до вподоби... Тільки мужам оцім не робіть нічого, бо на те вони прийшли під тінь даху мого.
GEN|19|9|А вони закричали: Іди собі геть! І сказали: Цей один був прийшов, щоб пожити чужинцем, а він став тут суддею! Тепер ми зло гірше тобі заподієм, ніж їм! І сильно вони налягали на мужа, на Лота, і підійшли, щоб висадити двері.
GEN|19|10|Тоді вистромили свою руку ті мужі, і впровадили Лота до себе до дому, а двері замкнули.
GEN|19|11|А людей, що при вході до дому зібрались, вони вдарили сліпотою, від малого аж до великого. І ті попомучилися, шукаючи входу.
GEN|19|12|І сказали ті мужі до Лота: Ще хто в тебе тут? Зятів і синів своїх, і дочок своїх, і все, що в місті твоє, виведи з цього місця,
GEN|19|13|бо ми знищимо це місце, бо збільшився їхній крик перед Господом, і Господь послав нас, щоб знищити його.
GEN|19|14|І вийшов Лот, і промовив до зятів своїх, що мали взяти дочок його, і сказав: Уставайте, вийдіть із цього місця, бо Господь знищить місто. Але в очах зятів він здавався як жартун.
GEN|19|15|А коли зійшла світова зірниця, то Анголи принагляли Лота, говорячи: Уставай, візьми жінку свою та обох дочок своїх, що знаходяться тут, щоб тобі не загинути через гріх цього міста.
GEN|19|16|А що він вагався, то ті мужі через Господню до нього любов схопили за руку його, і за руку жінки його, і за руку обох дочок його, і вивели його, і поставили поза містом.
GEN|19|17|І сталося, коли один з них виводив їх поза місто, то промовив: Рятуй свою душу, не оглядайся позад себе, і не затримуйся ніде в околиці. Ховайся на гору, щоб тобі не загинути.
GEN|19|18|А Лот їм відказав: Ні ж бо, Господи!
GEN|19|19|Ось Твій раб знайшов милість в очах Твоїх, і Ти побільшив Свою милість, що зробив її зо мною, щоб зберегти при житті мою душу; але я не встигну сховатись на гору, щоб бува не спіткало мене зло, і я помру.
GEN|19|20|Ось місто це близьке, щоб утекти туди, а воно маленьке. Нехай сховаюсь я туди, чи ж воно не маленьке? і буде жити душа моя.
GEN|19|21|І відказав Він до нього: Ось Я прихиливсь до твого прохання, щоб не зруйнувати міста, про яке ти казав.
GEN|19|22|Швидко сховайся туди, бо Я не зможу нічого зробити, аж поки не прийдеш туди. Тому й назвав ім'я тому місту: Цоар.
GEN|19|23|Сонце зійшло над землею, а Лот прибув до Цоару.
GEN|19|24|І Господь послав на Содом та Гомору дощ із сірки й огню, від Господа з неба.
GEN|19|25|І поруйнував ті міста, і всю околицю, і всіх мешканців міст, і рослинність землі.
GEN|19|26|А жінка його, Лотова, озирнулася позад нього, і стала стовпом соляним!...
GEN|19|27|І встав Авраам рано вранці, і подався до місця, де стояв був він перед лицем Господнім.
GEN|19|28|І він подивився на Содом та Гомору, і на всю поверхню землі тієї околиці. І побачив: ось здіймається дим від землі, немов дим із вапнярки...
GEN|19|29|І сталося, як нищив Бог міста тієї околиці, то згадав Бог Авраама, і вислав Лота з середини руїни, коли руйнував ті міста, що сидів у них Лот.
GEN|19|30|І піднявся Лот із Цоару, і осів на горі, й обидві дочки його з ним, бо боявся пробувати в Цоарі. І осів у печері, він та обидві дочки його.
GEN|19|31|І промовила старша молодшій: Наш батько старий, а чоловіка немає в цім краї, щоб прийшов до нас, як звичайно на цілій землі.
GEN|19|32|Ходи, напіймо свого батька вином, і покладімося з ним. І оживимо нащадків від нашого батька.
GEN|19|33|І ночі тієї вони напоїли вином свого батька. І прийшла старша та й поклалася з батьком своїм. А він не знав, коли вона лягла й коли встала...
GEN|19|34|І сталося другого дня, і старша сказала молодшій: Ось я минулої ночі поклалась була з своїм батьком. Напіймо його вином також ночі цієї, і прийди ти, покладися з ним, і оживимо нащадків від нашого батька.
GEN|19|35|І також ночі тієї вони напоїли вином свого батька. І встала молодша та й поклалася з ним. А він не знав, коли вона лягла й коли встала...
GEN|19|36|І завагітніли обидві Лотові дочки від батька свого.
GEN|19|37|І вродила старша сина, і назвала ім'я йому: Моав. Він батько моавів аж до цього дня.
GEN|19|38|А молодша вона вродила також, і назвала ймення йому: Бен-Аммі. Він батько синів Аммону аж до цього дня.
GEN|20|1|І вирушив звідти Авраам до краю Неґев поміж Кадешем і поміж Шуром, і оселився часово в Ґерарі.
GEN|20|2|І сказав Авраам на Сарру, жінку свою: Вона сестра моя. І послав Авімелех, цар Ґерару, і взяв Сарру.
GEN|20|3|І прийшов Бог до Авімелеха у сні нічнім, і сказав до нього: Ось ти вмираєш через жінку, яку взяв, бо вона має чоловіка.
GEN|20|4|А Авімелех не зближався до неї, і сказав: Господи, чи Ти вб'єш також люд праведний?
GEN|20|5|Чи ж не він був сказав мені: Вона моя сестра, а вона також вона сказала: Він мій брат. Я те зробив у невинності серця свого й у чистоті рук своїх.
GEN|20|6|І промовив до нього Бог у сні: І Я знаю, що в чистоті свого серця вчинив ти оце, і Я теж удержав тебе, щоб не згрішив проти Мене. Тому то не дав Я тобі доторкнутись до неї.
GEN|20|7|А тепер верни жінку цього мужа, бо він пророк, і буде молитися за тебе, і живи. А коли ти не вернеш, то знай, що справді помреш ти й усе, що твоє.
GEN|20|8|І встав Авімелех рано вранці, і покликав усіх рабів своїх, та й сказав усі ці слова до їхніх ушей. А люди ті сильно злякалися.
GEN|20|9|І закликав Авімелех Авраама, і промовив до нього: Що ти нам учинив? І чим згрішив я проти тебе, що ти приніс на мене й на царство моє великий гріх? Учинки, яких не роблять, ти зо мною вчинив!
GEN|20|10|І сказав Авімелех Авраамові: Що ти мав на увазі, що вчинив таку річ?
GEN|20|11|І сказав Авраам: Бо подумав я: Нема ж страху Божого в місцевості цій, тому вб'ють мене за жінку мою.
GEN|20|12|І притім вона справді сестра моя, вона дочка батька мого, тільки не дочка матері моєї, і стала за жінку мені.
GEN|20|13|І сталося, коли Бог учинив мене мандрівником з дому батька мого, то сказав я до неї: То буде твоя ласка, яку вчиниш зо мною: у кожній місцевості, куди прийдем, говори ти на мене: він мій брат.
GEN|20|14|І взяв Авімелех дрібну та велику худобу, і рабів та невільниць, та й дав Авраамові. І вернув йому Сарру, жінку його.
GEN|20|15|І сказав Авімелех: Ось край мій перед обличчям твоїм, осядь там, де тобі до вподоби.
GEN|20|16|А Саррі сказав: Ось тисячу секлів срібла я дав братові твоєму. Оце тобі накриття на очі перед усіма, хто з тобою. І перед усіма ти оправдана.
GEN|20|17|І помолився Авраам Богові, і вздоровив Бог Авімелеха, і жінку його, і невільниць його, і почали вони знову роджати.
GEN|20|18|Бо справді стримав був Господь кожну утробу Авімелехового дому через Сарру, Авраамову жінку.
GEN|21|1|А Господь згадав Сарру, як сказав був, і вчинив Господь Саррі, як Він говорив.
GEN|21|2|І Сарра зачала, і породила сина Авраамові в старості його на означений час, що про нього сказав йому Бог.
GEN|21|3|І назвав Авраам ім'я синові своєму, що вродився йому, що Сарра йому породила: Ісак.
GEN|21|4|І обрізав Авраам Ісака, сина свого, коли мав він вісім день, як Бог наказав був йому.
GEN|21|5|А Авраам був віку ста літ, як уродився йому Ісак, син його.
GEN|21|6|І промовила Сарра: Сміх учинив мені Бог, кожен, хто почує, буде сміятися з мене.
GEN|21|7|І промовила: Хто б сказав Авраамові: Сарра годує синів? Бо вродила я сина в старості його.
GEN|21|8|І дитина росла, і була відлучена. І справив Авраам велику гостину в день відлучення Ісака.
GEN|21|9|І побачила Сарра сина Аґари єгиптянки, що вродила була Авраамові, що він насміхається.
GEN|21|10|І сказала вона Авраамові: Прожени ту невільницю та сина її, бо не буде наслідувати син тієї невільниці разом із сином моїм, із Ісаком.
GEN|21|11|Але ця справа була дуже не до вподоби Авраамові через сина його.
GEN|21|12|І промовив Господь Авраамові: Нехай не буде не до вподоби тобі це через хлопця та через невільницю твою. Усе, що скаже тобі Сарра, послухай голосу її, бо Ісаком буде покликане тобі потомство.
GEN|21|13|І також сина невільниці тієї учиню його народом, бо він твоє насіння.
GEN|21|14|І встав рано Авраам, і взяв хліба й бурдюка води, і дав до Аґари на плече її, також дитину, та й послав її. І пішла вона, та й заблудила в пустині Беер-Шева.
GEN|21|15|І скінчилась вода в бурдюці, і покинула вона дитину під одним із кущів.
GEN|21|16|І пішла вона, і сіла собі навпроти, на віддалі як стрілити луком, бо сказала: Нехай я не бачу смерти цієї дитини! І сіла навпроти, і піднесла свій голос та й заплакала.
GEN|21|17|І почув Бог голос того хлопця. І кликнув до Аґари Божий Ангол із неба, і сказав їй: Що тобі, Аґаро? Не бійс, бо почув Бог голос хлопц, де він там.
GEN|21|18|Устань, підійми хлопця, і рукою своєю держи його, бо великим народом зроблю Я його.
GEN|21|19|І відкрив Бог очі її, і вона побачила криницю води. І пішла вона, і наповнила бурдюка водою, та й напоїла хлопця.
GEN|21|20|І з хлопцем був Бог, і він виріс. І осів у пустині, і став він стрілець-лучник.
GEN|21|21|І осів він у пустині Паран, а мати його взяла йому жінку з єгипетського краю.
GEN|21|22|І сталося часу того, і сказав Авімелех і Піхол, головний провідник його війська, до Авраама, говорячи: Бог із тобою в усьому, що ти робиш!
GEN|21|23|А тепер присягни ж мені Богом отут, що ти не обманиш мене, і нащадка мого, і онука мого. І яка була ласка, яку я до тебе чинив, ти вчиниш зо мною та з краєм, що ти в нім чужинцем пробуваєш.
GEN|21|24|І сказав Авраам: Я присягаю!
GEN|21|25|І Авраам дорікав Авімелехові за криницю води, що її відняли були Авімелехові раби.
GEN|21|26|І сказав Авімелех: Я не знаю, хто вчинив оту річ, ані ти не розповів мені, й ані я не чув, хібащо сьогодні.
GEN|21|27|І взяв Авраам дрібну та велику худобу, та й дав Авімелехові, і обидва вони склали умову.
GEN|21|28|І поставив Авраам сім овечок з дрібного товару осібно.
GEN|21|29|І сказав Авімелех до Авраама: Що вони, сім овечок отих, що ти їх поставив осібно?
GEN|21|30|А той відказав: Бо з моєї руки сім овечок ти візьмеш, щоб для мене були на свідоцтво, що я викопав цю криницю.
GEN|21|31|Тому то назвав він це місце Беер-Шева, бо там поклялися вони.
GEN|21|32|І склали умову вони в Беер-Шеві. І встав Авімелех та Піхол, головний провідник його війська, і вернулись вони до краю филистимського.
GEN|21|33|А Авраам посадив тамариска в Беер-Шеві, і кликав там Ім'я Господа, Бога Вічного.
GEN|21|34|І Авраам пробував у филистимській землі багато днів.
GEN|22|1|І сталось після цих випадків, що Бог випробовував Авраама. І сказав Він до нього: Аврааме! А той відказав: Ось я!
GEN|22|2|І промовив Господь: Візьми свого сина, свого одинака, що його полюбив ти, Ісака, та й піди собі до краю Морія, і принеси там його в цілопалення на одній із тих гір, що про неї скажу тобі.
GEN|22|3|І встав Авраам рано вранці, і свого осла осідлав; і взяв із собою двох слуг та Ісака, сина свого, і для цілопалення дров нарубав. І встав, і пішов він до місця, що про нього сказав йому Бог.
GEN|22|4|А третього дня Авраам звів очі свої, та й побачив те місце здалека.
GEN|22|5|І сказав Авраам своїм слугам: Сідайте собі тут з ослом, а я й хлопець підем аж туди, і поклонимося, і повернемося до вас.
GEN|22|6|І взяв Авраам дрова для цілопалення, і поклав на Ісака, сина свого, і взяв в свою руку огонь та ножа, і пішли вони разом обоє.
GEN|22|7|І сказав Ісак до Авраама, свого батька, говорячи: Батьку мій! А той відказав: Ось я, сину мій! І промовив Ісак: Ось огонь та дрова, а де ж ягня на цілопалення?
GEN|22|8|І відказав Авраам: Бог нагледить ягня Собі на цілопалення, сину мій! І пішли вони разом обоє.
GEN|22|9|І вони прийшли до місця, що про нього сказав йому Бог. І збудував там Авраам жертівника, і дрова розклав, і зв'язав Ісака, сина свого, і поклав його на жертівника над дровами.
GEN|22|10|І простяг Авраам свою руку, і взяв ножа, щоб зарізати сина свого...
GEN|22|11|Та озвався до нього Ангол Господній із неба й сказав: Аврааме, Аврааме! А той відізвався: Ось я!
GEN|22|12|І Ангол промовив: Не витягай своєї руки до хлопця, і нічого йому не чини, бо тепер Я довідався, що ти богобійний, і не пожалів для Мене сина свого, одинака свого.
GEN|22|13|А Авраам звів очі свої та й побачив, аж ось один баран зав'яз у гущавині своїми рогами. І пішов Авраам, і взяв барана, і приніс його на цілопалення замість сина свого.
GEN|22|14|І назвав Авраам ім'я місця того: Господь нагледить, що й сьогодні говориться: На горі Господь з'явиться.
GEN|22|15|А Ангол Господній із неба озвався до Авраама подруге,
GEN|22|16|і сказав: Клянуся Собою, це слово Господнє, тому, що вчинив ти цю річ, і не пожалів був сина свого, одинака свого,
GEN|22|17|то благословляючи, Я поблагословлю тебе, і розмножуючи, розмножу потомство твоє, немов зорі на небі, і немов той пісок, що на березі моря. І потомство твоє внаслідує брами твоїх ворогів.
GEN|22|18|І всі народи землі будуть потомством твоїм благословляти себе через те, що послухався ти Мого голосу.
GEN|22|19|І вернувсь Авраам до слуг своїх.
GEN|22|20|І сталося по тих випадках, і сказано Авраамові так: Ось також Мілка вродила синів Нахорові, братові твоєму:
GEN|22|21|Уца, перворідного його, і Буза, брата його, і Кемуїла, батька Арамового,
GEN|22|22|І Кеседа, і Хазо, і Пілдаша, і Їдлафа, і Бетуїла.
GEN|22|23|А Бетуїл породив Ревеку. Цих восьмерох породила Мілка Нахорові, братові Авраамовому.
GEN|22|24|А наложниця його а їй на ймення Реума вродила й вона Теваха й Ґахама, і Тахаша й Мааху.
GEN|23|1|І було життя Сарриного сто літ і двадцять літ і сім літ, літа життя Сарриного.
GEN|23|2|І вмерла Сарра в Кіріят-Арбі, це Хеврон у Краї ханаанському. І прибув Авраам голосити над Саррою та плакати за нею.
GEN|23|3|І встав Авраам від обличчя небіжки своєї, та й сказав синам Хетовим, говорячи:
GEN|23|4|Я приходько й захожий між вами. Дайте в себе мені власність для гробу, і нехай я поховаю свою небіжку з-перед обличчя свого.
GEN|23|5|І відповіли сини Хетові Авраамові, та й сказали йому:
GEN|23|6|Послухай нас, пане мій, ти Божий князь серед нас! У добірнім із наших гробів поховай небіжку свою. Ніхто з нас не затримає гробу свого від тебе, щоб поховати небіжку твою.
GEN|23|7|І встав Авраам, і вклонився народу тієї землі, синам Хетовим,
GEN|23|8|та й промовив до них і сказав: Коли ви згідні поховати небіжку мою з-перед обличчя мого, то послухайте мене, і настирливо просіть для мене Ефрона, сина Цохарового,
GEN|23|9|і нехай мені дасть він печеру Махпелу, що його, що в кінці його поля, за гроші повної ваги, хай мені її дасть поміж вами на власність для гробу.
GEN|23|10|А Ефрон пробував серед Хетових синів. І відповів хіттеянин Ефрон Авраамові, так що чули сини Хетові й усі, хто входив у браму його міста, говорячи:
GEN|23|11|Ні, пане мій, послухай мене! Поле віддав я тобі, і печеру, що на нім, віддав я тобі, на очах синів народу мого я віддав її тобі. Поховай небіжку свою.
GEN|23|12|І вклонивсь Авраам перед народом тієї землі,
GEN|23|13|та й сказав до Ефрона, так що чув був народ тієї землі, говорячи: Коли б тільки мене ти послухав! Я дам срібло за поле, візьми ти від мене, і хай поховаю небіжку свою.
GEN|23|14|А Ефрон відповів Авраамові, говорячи йому:
GEN|23|15|Пане мій, послухай мене! Земля чотирьох сотень шеклів срібла, що вона поміж мною та поміж тобою? А небіжку свою поховай!
GEN|23|16|І послухав Авраам Ефрона. І відважив Авраам Ефронові срібло, про яке той був сказав, так що чули сини Хетові, чотири сотні шеклів срібла купецької ваги.
GEN|23|17|І стало поле Ефронове, що в Махпелі воно, що перед Мамре, поле й печера, що на ньому, і кожне дерево, що в полі, що в усій границі його навколо,
GEN|23|18|купном Авраамові в присутності синів Хетових, усіх, хто входив до брами міста його.
GEN|23|19|І по цьому Авраам поховав Сарру, жінку свою, в печері поля Махпели, перед Мамре, це Хеврон у землі ханаанській.
GEN|23|20|І стало поле й печера, що на нім, Авраамові на власність для гробу від синів Хетових.
GEN|24|1|А Авраам був старий, у літа ввійшов. І Господь Авраама поблагословив був усім.
GEN|24|2|І сказав Авраам до свого раба, найстаршого дому свого, що рядив над усім, що він мав: Поклади свою руку під стегно моє,
GEN|24|3|і я заприсягну тебе Господом, Богом неба й Богом землі, що ти не візьмеш жінки для сина мого з-посеред дочок ханаанеянина, серед якого я пробуваю.
GEN|24|4|Бо ти підеш до краю мого, і до місця мого народження, і візьмеш жінку для сина мого, для Ісака.
GEN|24|5|І сказав раб до нього: Може та жінка не схоче за мною піти до цієї землі, то чи справді поверну я твого сина до краю, звідки ти вийшов?
GEN|24|6|І промовив до нього Авраам: Стережися, щоб ти не вернув мого сина туди!
GEN|24|7|Господь, що взяв мене з дому батька мого й з краю мого народження, і що промовляв був до мене, і що присягнув мені, кажучи: Твоїм нащадкам Я дам оцю землю, Він пошле Свого Ангола перед обличчям твоїм, і ти візьмеш звідти жінку для сина мого!
GEN|24|8|А коли ота жінка не схоче піти за тобою, то ти будеш очищений з цієї присяги своєї. Тільки сина мого ти туди не вертай.
GEN|24|9|І раб поклав свою руку під стегно Авраама, пана свого, і йому присягнув на цю справу.
GEN|24|10|І взяв той раб десять верблюдів із верблюдів пана свого, та й пішов. І взяв різне добро свого пана в руку свою. І він устав, і пішов в Месопотамію до міста Нахора.
GEN|24|11|І поставив верблюди навколішки за містом при водній криниці надвечір, на час, як виходять жінки воду брати,
GEN|24|12|та й промовив: Господи, Боже пана мого Авраама, подай же сьогодні мені це, і милість вчини з паном моїм Авраамом!
GEN|24|13|Ось я стою над водним джерелом, а дочки мешканців міста виходять воду брати.
GEN|24|14|І станеться, що дівчина, до якої скажу: Нахили но глека свого, я нап'юся, а вона відповість: Пий, і так само верблюди твої я понапуваю, її Ти призначив для раба Свого, для Ісака. І з цього пізнаю, що Ти милість учинив з моїм паном.
GEN|24|15|І сталося, поки він закінчив говорити, аж ось виходить Ревека, що була народжена Бетуїлові, синові Мілки, жінки Нахора, Авраамового брата. А її глек на плечі в неї.
GEN|24|16|А дівчина та вельми вродлива з обличчя; була дівиця, і чоловік не пізнав ще її. І зійшла вона до джерела, і наповнила глека свого, та й вийшла.
GEN|24|17|І вибіг той раб назустріч їй, та й сказав: Дай но напитись води з твого глека!
GEN|24|18|А та відказала: Напийся, мій пане! І вона поспішила, і зняла свого глека на руку свою, і напоїла його.
GEN|24|19|А коли закінчила поїти його, то сказала: Також для верблюдів твоїх наберу я води, аж поки вони не нап'ються.
GEN|24|20|І метнулась вона, і глека свого спорожнила до пійла. І ще до криниці побігла набрати, і набрала води всім верблюдам його.
GEN|24|21|А чоловік той дивувався їй та мовчав, щоб пізнати, чи Господь пощастив дорогу йому, чи ні?
GEN|24|22|І сталося, як перестали верблюди пити, то взяв той чоловік золоту сережку, пів шекля вага їй, і два наручні на руки її, на десять шеклів золота вага їм,
GEN|24|23|та й сказав: Чия ти дочка? Скажи ж мені, чи в домі батька твойого є місце для нас ночувати?
GEN|24|24|Вона відказала йому: Я дочка Бетуїла, сина Мілки, що його породила вона для Нахора.
GEN|24|25|І сказала до нього: І соломи, і паші багато є в нас, також місце ночувати.
GEN|24|26|І той чоловік нахилився, і вклонився Богові аж до землі,
GEN|24|27|та й сказав: Благословенний Господь, Бог пана мого Авраама, що не опустив милости Своєї й вірности Своєї від пана мого! Я був у дорозі, Господь припровадив мене до дому братів мого пана.
GEN|24|28|І побігла дівчина, і розповіла в домі своєї матері про цю пригоду.
GEN|24|29|А в Ревеки був брат, на ймення йому Лаван. І побіг Лаван до того чоловіка надвір, до джерела.
GEN|24|30|І сталося, як він побачив сережку та наручні на руках сестри своєї, і коли почув слова Ревеки, сестри своєї, що говорила: Отак говорив мені той чоловік, то прибув він до того чоловіка, а той ось стоїть при верблюдах біля джерела,
GEN|24|31|і сказав: Увійди, благословенний Господа! Чого стоятимеш надворі? А я опорожнив дім і місце для верблюдів.
GEN|24|32|І ввійшов той чоловік до дому. А Лаван порозсідлував верблюди, і дав соломи й паші для верблюдів, і води, щоб умити ноги йому й ноги людям, що були з ним.
GEN|24|33|І поставлено перед ним, щоб він їв. А той відказав: Не буду їсти, аж поки не розкажу своєї справи. А Лаван відказав: Говори!
GEN|24|34|І той став говорити: Я раб Авраамів.
GEN|24|35|А Господь щедро поблагословив мого пана, і він став великий. І дав Він йому худобу дрібну та велику, і срібло, і золото, і рабів, і невільниць, і верблюди, й осли.
GEN|24|36|А Сарра, жінка пана мого, бувши старою, уродила панові моєму сина. А він йому все дав, що мав.
GEN|24|37|І заприсяг мене пан мій, говорячи: Не візьмеш жінки для сина мого з-посеред дочок ханаанеянина, що я пробуваю в його краю.
GEN|24|38|Але підеш до дому батька мого, і до мого роду, і візьмеш жінку для сина мого.
GEN|24|39|І сказав я до пана свого: Може та жінка не піде за мною?
GEN|24|40|І сказав він до мене: Господь, що ходив перед обличчям моїм, пошле Свого Ангола з тобою, і дорогу твою пощастить, і ти візьмеш жінку для сина мого з роду мого й з дому батька мого.
GEN|24|41|Тоді будеш очищений ти від закляття мого, як прийдеш до роду мого, а коли вони не дадуть тобі, то будеш ти чистий від закляття мого.
GEN|24|42|І прибув я сьогодні до джерела, та й сказав: Господи, Боже пана мого Авраама, коли б же Ти вчинив щасливою дорогу мою, що нею ходжу я!
GEN|24|43|Ось я стою над джерелом води, і станеться, що дівчина, яка вийде води брати, а я їй скажу: Дай но мені напитися трохи води з свого глека,
GEN|24|44|вона ж відкаже мені: Пий і ти, і для верблюдів твоїх наберу я води, то вона та жінка, яку призначив Господь для сина пана мого.
GEN|24|45|І поки скінчив я говорити в своїм серці, аж ось виходить Ревека, а її глек на плечі в неї. І зійшла вона до джерела, та й набрала води. І сказав я до неї: Напій же мене!
GEN|24|46|І метнулась вона, і свого глека з себе зняла та й сказала: Пий, а я понапуваю й верблюди твої. І я пив, а вона понапувала й ті верблюди.
GEN|24|47|А я запитався її та й сказав: Чия ти дочка? А вона відказала: Я дочка Бетуїла, сина Нахорового, якого породила йому Мілка. І сережку надів я до носа її, і наручні на руки її.
GEN|24|48|І я нахилився, і вклонився до землі Господеві, і поблагословив Господа, Бога пана мого Авраама, що Він провадив мене дорогою визначеною, щоб узяти дочку брата пана мого для сина його.
GEN|24|49|А тепер, якщо милосердя та правду ви чините з паном моїм, то скажіть мені; коли ж ні, то скажіть мені, і я звернуся праворуч або ліворуч.
GEN|24|50|І відповіли Лаван і Бетуїл та й сказали: Від Господа вийшла та річ, ми не можем сказати тобі нічого злого чи доброго.
GEN|24|51|Ось перед тобою Ревека, візьми та й іди, і нехай вона стане за жінку синові пана твого, як Господь говорив був.
GEN|24|52|І сталося, коли їхні слова почув раб Авраамів, то вклонивсь до землі Господеві.
GEN|24|53|І вийняв той раб срібний посуд, і посуд золотий та шати, і дав Ревеці, і дав цінні речі братові її та матері її.
GEN|24|54|І їли й пили він та люди, що з ним, і ночували. А коли рано встали, то він сказав: Відішліть мене до пана мого.
GEN|24|55|І сказав її брат та мати її: Нехай посидить дівчина з нами хоч днів з десять, потім підеш.
GEN|24|56|І сказав він до них: Не спізняйте мене, бо Господь пощастив мою путь. Відішліть мене, і нехай я піду до пана свого.
GEN|24|57|А вони відказали: Покличмо дівчину, і запитаймо її саму.
GEN|24|58|І покликали Ревеку, і сказали до неї: Чи ти підеш з оцим чоловіком? А вона відказала: Піду.
GEN|24|59|І послали вони Ревеку, сестру свою, і няньку її, і раба Авраамового, і людей його.
GEN|24|60|І вони поблагословили Ревеку й сказали до неї: Ти наша сестра, будь матір'ю для тисячі десятків тисяч, і нехай нащадки твої внаслідують брами твоїх ворогів.
GEN|24|61|І встала Ревека й служниці її, і посідали на верблюдів, і поїхала за тим чоловіком. І взяв раб Ревеку й відійшов.
GEN|24|62|А Ісак був вернувся з подорожі до криниці Лахай-Рої, і сидів у краї південному.
GEN|24|63|І вийшов Ісак на прогулянку в поле, як вечір наставав. І він звів свої очі, і побачив, ось верблюди йдуть.
GEN|24|64|І Ревека звела свої очі, та й Ісака побачила, і злізла з верблюда.
GEN|24|65|І сказала вона до раба: Хто отой чоловік, що полем іде нам назустріч? А раб відповів: То мій пан. І вона покривало взяла, та й накрилась.
GEN|24|66|І раб розповів Ісакові про всі речі, які він учинив.
GEN|24|67|І впровадив її Ісак до намету Сарри, матері своєї. І взяв він Ревеку, і за жінку йому вона стала, і він її покохав. І Ісак був утішений по смерті матері своєї.
GEN|25|1|А Авраам іще взяв жінку, а ймення їй Кетура.
GEN|25|2|А вона породила йому Зімрана, і Йокшана, і Мадана, і Мідіяна, і Їшбака, і Шуаха.
GEN|25|3|А Йокшан породив був Шеву та Дедана. А сини Деданові були: ашшури, і летуші, і леуми.
GEN|25|4|А сини Мідіянові: Ефа, і Ефер, і Ханох, і Авіда, і Елдаа, усі вони сини Кетури.
GEN|25|5|І віддав Авраам усе, що мав, Ісакові.
GEN|25|6|А синам наложниць, що були в Авраама, дав Авраам подарунки, і відіслав їх від Ісака, сина свого, коли сам ще живий був, на схід, до краю східнього.
GEN|25|7|А оце дні літ Авраамового життя, які він прожив: сто літ, і сімдесят літ, і п'ять літ.
GEN|25|8|І спочив та й умер Авраам у старощах добрих, старий і нажившись. І він прилучився до своєї рідні.
GEN|25|9|І поховали його Ісак та Ізмаїл, сини його, у печері Махпелі, на полі Ефрона, сина Цохара хіттеянина, що навпроти Мамре,
GEN|25|10|поле, що його Авраам був купив від синів Хетових, там був похований Авраам і Сарра, жінка його.
GEN|25|11|І сталося по Авраамовій смерті, і поблагословив Бог Ісака, сина його. І осів Ісак при криниці Лахай-Рої.
GEN|25|12|А оце нащадки Ізмаїла, Авраамового сина, що його породила Авраамові єгиптянка Аґар, невільниця Саррина.
GEN|25|13|І оце імена синів Ізмаїла, за їхніми іменами й за нащадками їх: перворідний Ізмаїлів Невайот, і Кедар, і Адбеїл, і Мівсам,
GEN|25|14|І Мішма, і Дума, і Масса,
GEN|25|15|Хадад, і Тема, Єтур, Нафіш, і Кедма.
GEN|25|16|Оце вони, сини Ізмаїлові, і їхні ймення за дворами їх і за їх кочовищами, дванадцять начальників для їхніх племен.
GEN|25|17|А оце літа життя Ізмаїлового: сто літ, і тридцять літ, і сім літ. І спочив та й умер він, і був узятий до своєї рідні.
GEN|25|18|І розложилися вони від Хавіли аж до Шуру, що навпроти Єгипту, як іти до Ашшуру. І він оселився перед усіма своїми братами.
GEN|25|19|А оце оповість про Ісака, Авраамового сина. Авраам породив Ісака.
GEN|25|20|І був Ісак віку сорока літ, як він узяв собі за жінку Ревеку, дочку Бетуїла арамеянина, з Падану арамейського, сестру арамеянина Лавана.
GEN|25|21|І молився Ісак до Господа про жінку свою, бо неплідна була. І Господь був ублаганий ним, і завагітніла Ревека, жінка його.
GEN|25|22|І кидалися діти в утробі її. І сказала вона: Коли так, то для чого я це переношу? І пішла запитатися Господа.
GEN|25|23|І промовив до неї Господь: Два племена в утробі твоїй, і два народи з твого нутра будуть виділені, і стане сильніший народ від народу, і старший молодшому буде служити.
GEN|25|24|І сповнились дні її, щоб родити, і ось близнюки в утробі її.
GEN|25|25|І вийшов перший червонуватий, увесь він немов плащ волосяний. І назвали ймення йому: Ісав.
GEN|25|26|А потім вийшов його брат, а рука його трималася п'яти Ісава. І назвав ім'я йому: Яків. А Ісак був віку шостидесяти літ, коли народились вони.
GEN|25|27|І виросли хлопці. І став Ісав чоловіком, що знався на вловах, чоловіком поля, а Яків чоловіком мирним, що в наметах сидів.
GEN|25|28|І полюбив Ісак Ісава, бо здобич мисливська його йому смакувала, а Ревека любила Якова.
GEN|25|29|І зварив був Ісак їжу, а з поля прибув Ісав, і змучений був.
GEN|25|30|І сказав Ісав до Якова: Нагодуй мене отим червоним, червоним отим, бо змучений я. Тому то назвали ймення йому: Едом.
GEN|25|31|А Яків сказав: Продай же нині мені своє перворідство.
GEN|25|32|І промовив Ісав: Ось я умираю, то нащо ж мені оте перворідство?
GEN|25|33|А Яків сказав: Присягни ж мені нині. І той присягнув йому, і продав перворідство своє Якову.
GEN|25|34|І Яків дав Ісавові хліба й сочевичного варива. А той з'їв, і випив, і встав та й пішов. І знехтував Ісав перворідство своє.
GEN|26|1|І настав був голод у Краю, окрім голоду першого, що був за днів Авраамових. І пішов Ісак до Авімелеха, царя филистимського, до Ґерару.
GEN|26|2|І явився йому Господь і сказав: Не ходи до Єгипту, оселися в землі, про яку Я скажу тобі.
GEN|26|3|Оселися хвилево в землі тій, і Я буду з тобою, і тебе поблагословлю, бо тобі та нащадкам твоїм дам усі оці землі. І Я виконаю присягу, що нею поклявся був Авраамові, батьку твоєму.
GEN|26|4|І розмножу нащадків твоїх, немов зорі на небі, і потомству твоєму Я дам усі оці землі. І поблагословляться в потомстві твоїм усі народи землі,
GEN|26|5|через те, що Авраам послухав Мого голосу, і виконував те, що виконувати Я звелів: заповіді Мої, постанови й закони Мої.
GEN|26|6|І осів Ісак у Ґерарі.
GEN|26|7|І питалися люди тієї місцевости про жінку його. А він відказав: Вона сестра моя, бо боявся сказати: Вона жінка моя, щоб не вбили мене люди тієї місцевости через Ревеку, бо вродлива з обличчя вона.
GEN|26|8|І сталося, коли він там довго жив, і дивився Авімелех, цар филистимський, через вікно, та й побачив, ось Ісак забавляється з Ревекою, жінкою своєю.
GEN|26|9|І покликав Авімелех Ісака та й сказав: Тож оце вона жінка твоя! А як ти сказав був: Вона сестра моя? Ісак же йому відповів: Бо сказав, щоб не вмерти мені через неї!
GEN|26|10|І сказав Авімелех: Що ж то нам учинив ти? Один із народу був мало не ліг із твоєю жінкою, і ти гріх би спровадив на нас!
GEN|26|11|І наказав Авімелех усьому народові, говорячи: Хто доторкнеться цього чоловіка та жінки його, той певно буде забитий.
GEN|26|12|І посіяв Ісак у землі тій, і зібрав того року стокротно, і Господь поблагословив був його.
GEN|26|13|І забагатів оцей чоловік, і багатів усе більше, аж поки не став сильно багатий.
GEN|26|14|І була в нього отара овець та кіз, і череда товару, і багато рабів. І заздрили йому филистимляни.
GEN|26|15|І всі криниці, що їх повикопували раби батька його, за днів батька його Авраама, филистимляни позатикали, і понаповнювали їх землею.
GEN|26|16|І сказав Авімелех Ісакові: Іди ти від нас, бо зробився ти значно сильніший за нас!
GEN|26|17|І пішов Ісак звідти, і в долині Ґерару розтаборився, та й осів там.
GEN|26|18|І знову Ісак повикопував криниці на воду, що їх повикопували були за днів батька його Авраама, а позатикали були їх филистимляни по Авраамовій смерті. І він назвав їм імення, як імення, що батько його був їм назвав.
GEN|26|19|І копали Ісакові раби в долині, і знайшли там криницю живої води.
GEN|26|20|І сварилися пастухи ґерарські з пастухами Ісаковими, кажучи: Це наша вода! І він назвав ім'я для тієї криниці: Есек, бо сварилися з ним.
GEN|26|21|І викопали вони іншу криницю, і сварилися також за неї. І він назвав для неї ім'я: Ситна.
GEN|26|22|І він пересунувся звідти, і викопав іншу криницю, і не сварились за неї. І він назвав для неї ім'я: Реховот, і сказав: Тепер нам поширив Господь, і в Краю ми розмножимось.
GEN|26|23|А звідти піднявся він до Беер-Шеви.
GEN|26|24|І явився йому Господь тієї ночі й сказав: Я Бог Авраама, батька твого; не бійся, бо Я з тобою! І поблагословлю Я тебе, і розмножу нащадків твоїх ради Авраама, Мойого раба.
GEN|26|25|І він збудував там жертівника, і покликав Господнє Ймення. І поставив він там намета свого, а раби Ісакові криницю там викопали.
GEN|26|26|І прийшов до нього з Ґерару Авімелех, і Ахуззат, товариш його, і Піхол, головний начальник війська його.
GEN|26|27|І сказав їм Ісак: Чого ви до мене прийшли? Ви ж зненавиділи мене, і вислали мене від себе.
GEN|26|28|А ті відказали: Ми бачимо справді, що з тобою Господь. І ми сказали: Нехай буде клятва поміж нами, поміж нами й поміж тобою, і складімо умову з тобою,
GEN|26|29|що не вчиниш нам злого, як і ми не торкнулись до тебе, і як ми робили з тобою тільки добро, і тебе відіслали з миром. Ти тепер благословенний від Господа!
GEN|26|30|І він учинив для них гостину, і вони їли й пили.
GEN|26|31|А рано вони повставали, і присягли один одному. І відіслав їх Ісак, і вони пішли від нього з миром.
GEN|26|32|І сталося того дня, і прийшли Ісакові раби, і розказали йому про криницю, яку вони викопали. І сказали йому: Ми воду знайшли!
GEN|26|33|І він назвав її: Шів'а, чому ймення міста того Беер-Шева аж до сьогоднішнього дня.
GEN|26|34|І був Ісав віку сорока літ, і взяв жінку Єгудиту, дочку хіттеянина Беері, і Босмату, дочку хіттеянина Елона.
GEN|26|35|І вони стали гіркотою духа для Ісака й Ревеки.
GEN|27|1|І сталося, що зостарівсь Ісак, і затемнились очі йому, і він не бачив. І покликав він старшого сина свого Ісава, і промовив до нього: Мій сину! А той відказав йому: Ось я!
GEN|27|2|І промовив до нього Ісак: Оце я зостарівся, не знаю дня смерти своєї...
GEN|27|3|А тепер візьми знаряддя своє, сагайдака свого й лука свого, та й вийди на поле, і злови мені здобич мисливську.
GEN|27|4|І зготуй мені наїдок смачний, як я люблю, і принеси мені, і нехай я з'їм, щоб поблагословила тебе душа моя, поки помру.
GEN|27|5|А Ревека чула, як говорив Ісак до Ісава, сина свого. І пішов Ісав на поле, щоб зловити й принести здобич мисливську.
GEN|27|6|А Ревека сказала Якову, синові своєму, говорячи: Ось я чула, як твій батько казав до Ісава, брата твого, говорячи:
GEN|27|7|Принеси но здобич мисливську мені, і зроби мені наїдок смачний, нехай з'їм, і поблагословлю тебе перед лицем Господнім перед смертю своєю.
GEN|27|8|А тепер, сину мій, послухай мого голосу, те, що я розкажу тобі.
GEN|27|9|Іди до отари, і візьми мені звідти двоє добрих козлят, а я їх приготую, як наїдок смачний для батька твого, як він любить.
GEN|27|10|І принесеш батькові своєму, і буде він їсти, щоб поблагословити тебе перед смертю своєю.
GEN|27|11|І промовив Яків до Ревеки, матері своєї: Таж брат мій Ісав чоловік волохатий, а я чоловік гладенький!
GEN|27|12|Може обмацає мене батько мій, і я стану в очах його як обманець, і спроваджу на себе прокляття, а не благословення...
GEN|27|13|І сказала йому його мати: На мені прокляття твоє, сину мій! Тільки послухай слів моїх, та йди принеси мені.
GEN|27|14|І пішов він, і взяв, і приніс своїй матері. І зробила мати його наїдок смачний, як любив його батько.
GEN|27|15|І взяла Ревека гарні вбрання свого старшого сина Ісава, що були в домі з нею, і вбрала молодшого сина свого Якова.
GEN|27|16|А шкури козлят наділа на руки йому, і на гладеньку шию його.
GEN|27|17|І дала смачний наїдок та хліб, що вона спорядила, у руку Якова, сина свого.
GEN|27|18|І прибув він до батька свого та й сказав: Батьку мій! А той відказав: Ось я. Хто ти, мій сину?
GEN|27|19|А Яків промовив до батька свого: Я Ісав перворідний. Я зробив, як сказав ти мені. Уставай, сядь і попоїж із здобичі мисливської, щоб душа твоя поблагословила мене.
GEN|27|20|І сказав Ісак до сина свого: Як це ти так швидко знайшов, сину мій? А той відказав: Бо мені допоміг Господь, Бог твій.
GEN|27|21|І промовив Ісак до Якова: Підійди но, і нехай я обмацаю тебе, сину мій, чи ти це син мій Ісав, чи ні.
GEN|27|22|І підійшов Яків до Ісака, батька свого. А той обмацав його та й сказав: Голос голос Яковів, а руки руки Ісавові.
GEN|27|23|І не впізнав він його, бо були його руки як руки Ісава, брата його, волохаті, і поблагословив він його.
GEN|27|24|І сказав він: То ти син мій Ісав? А той відказав: Я.
GEN|27|25|І промовив Ісак: Подай же мені, і нехай з'їм з мисливської здобичі сина мого, щоб поблагословила тебе душа моя. І подав він йому, і він їв, і приніс йому вина, і він пив.
GEN|27|26|І промовив до нього Ісак, його батько: Підійди ж, і поцілуй мене, сину мій!
GEN|27|27|І він підійшов, і поцілував його. А той понюхав запах вбрання його, і поблагословив його, та й сказав: Дивись, запах сина мого немов запах поля, що його Господь благословив!
GEN|27|28|І хай Бог тобі дасть з роси Неба, і з ситости землі, і збіжжя багато й вина молодого!
GEN|27|29|Нехай тобі служать народи, і народи нехай тобі кланяються! Будь паном для братів своїх, і нехай тобі кланяються сини матері твоєї. Хто тебе проклинає проклятий, а хто поблагословить тебе благословенний!.
GEN|27|30|І сталося, як закінчив був Ісак благословляти Якова, і сталося, тільки но вийшов був Яків від обличчя Ісака, батька свого, аж Ісав, його брат, прийшов з полювання свого...
GEN|27|31|І також він приготовив наїдок смачний, і батьку своєму приніс. І сказав він до батька свого: Нехай встане мій батько, і хай їсть із здобичі мисливської сина свого, щоб душа твоя благословила мене!
GEN|27|32|І озвався до нього Ісак, його батько: Хто ти? А той відказав: Я син твій, твій перворідний Ісав.
GEN|27|33|І Ісак затремтів тремтінням аж надто великим, та й сказав: Хто ж тоді той, що мисливську здобич зловив, і до мене приніс, а я попоїв від усього, поки прийшов ти, і я поблагословив його? І він буде благословенний!
GEN|27|34|Як Ісав почув слова батька свого, то закричав криком сильним та вельми гірким. І сказав він до батька свого: Поблагослови мене, також мене, батьку мій!
GEN|27|35|А той відказав: Обманом прийшов був твій брат, та й забрав благословення твоє!
GEN|27|36|І промовив Ісав: Тому звалось ім'я його: Яків, і він обманив два рази мене: забрав перворідство моє, а це тепер забрав благословення моє. І сказав він: Чи ти не заховав для мене благословення?
GEN|27|37|А Ісак відповів і промовив до Ісава: Тож я вчинив його паном для тебе, та дав йому всіх братів його за рабів. І я забезпечив його хлібом і молодим вином. А що ж тоді тобі я зроблю, сину мій?
GEN|27|38|І сказав Ісав до батька свого: Чи в тебе одне те благословення, батьку мій? Поблагослови мене, також мене, батьку мій! І підніс Ісав голос свій, та й заплакав...
GEN|27|39|І відповів Ісак, батько його, та й промовив до нього: Ото буде садиба твоя без ситости землі, і без роси небесної згори.
GEN|27|40|І зо свого меча будеш жити, і будеш служити ти брату своєму. Та однако коли постараєшся, то зламаєш ярмо його з шиї своєї...
GEN|27|41|І зненавидів Ісав Якова через благословення, що поблагословив його батько його. І сказав Ісав у серці своєму: Нехай наближаться дні жалоби по батьку моєму, і я вб'ю Якова, брата свого.
GEN|27|42|І розказано Ревеці слова Ісава, її старшого сина. І послала, і покликала Якова, молодшого сина свого, та й сказала до нього: Ось Ісав, брат твій, тішиться тим, що уб'є тебе.
GEN|27|43|А тепер, сину мій, послухай мого голосу, і встань, і втечи собі до Лавана, брата мого, до Харану.
GEN|27|44|І посидиш у нього кілька часу, аж поки відвернеться лютість твого брата,
GEN|27|45|аж поки відвернеться гнів твого брата від тебе, і він забуде, що ти зробив був йому. Тоді я пошлю й заберу тебе звідти. Чого маю я стратити вас обох одного дня?
GEN|27|46|І сказала Ревека Ісакові: Життя мені обридло через дочок Хетових. Коли Яків візьме жінку з дочок Хетових, як ці, з дочок цього Краю, то нащо й жити мені?
GEN|28|1|І покликав Ісак Якова, і поблагословив його, і наказав йому та й промовив: Не бери жінки з дочок ханаанських.
GEN|28|2|Устань, піди до Падану арамейського, до дому Бетуїла, батька твоєї матері, і візьми собі звідти жінку з дочок Лавана, брата матері твоєї.
GEN|28|3|А Бог Всемогутній поблагословить тебе, і розплодить тебе, і розмножить тебе, і ти станеш громадою народів.
GEN|28|4|І дасть тобі благословення Авраамове, тобі та потомству твоєму з тобою, щоб віддати тобі землю твого тимчасового замешкання, що Бог дав був її Авраамові.
GEN|28|5|І послав Ісак Якова, і пішов він до Падану арамейського, до Лавана, сина Бетуїлового, арамеянина, брата Ревеки, матері Якова й Ісава.
GEN|28|6|І побачив Ісав, що Ісак поблагословив Якова, і послав його до Падану арамейського, щоб узяв собі звідти жінку, і поблагословив його, кажучи: Не бери жінки з дочок ханаанських,
GEN|28|7|і що послухався Яків батька свого й матері своєї, та й пішов до Падану арамейського.
GEN|28|8|І побачив Ісав, що дочки ханаанські недобрі в очах Ісака, батька його,
GEN|28|9|і пішов Ісав до Ізмаїла, і взяв Махалату, дочку Ізмаїла, сина Авраамового, сестру Невайотову, до жінок своїх за жінку.
GEN|28|10|І вийшов Яків із Беер-Шеви, і пішов до Харану.
GEN|28|11|І натрапив він був на одне місце, і ночував там, бо сонце зайшло було. І взяв він з каміння того місця, і поклав собі в голови. І він ліг на тім місці.
GEN|28|12|І снилось йому, ось драбина поставлена на землю, а верх її сягав аж неба. І ось Анголи Божі виходили й сходили по ній.
GEN|28|13|І ото Господь став на ній і промовив: Я Господь, Бог Авраама, батька твого, і Бог Ісака. Земля, на якій ти лежиш, Я дам її тобі та нащадкам твоїм.
GEN|28|14|І буде потомство твоє, немов порох землі. І поширишся ти на захід, і на схід, і на північ, і на південь. І благословляться в тобі та в нащадках твоїх всі племена землі.
GEN|28|15|І ось Я з тобою, і буду тебе пильнувати скрізь, куди підеш, і верну тебе до цієї землі, бо Я не покину тебе, аж поки не вчиню, що Я сказав був тобі.
GEN|28|16|І прокинувся Яків зо свого сну, та й сказав: Дійсно, Господь пробуває на цьому місці, а того я й не знав!
GEN|28|17|І злякався він і сказав: Яке страшне оце місце! Це ніщо інше, як дім Божий, і це брама небесна.
GEN|28|18|І встав Яків рано вранці, і взяв каменя, що поклав був собі в голови, і поставив його за пам'ятника, і вилив оливу на його верх.
GEN|28|19|І назвав він ім'я тому місцю: Бет-Ел, а ймення того міста напочатку було Луз.
GEN|28|20|І склав Яків обітницю, говорячи: Коли Бог буде зо мною, і буде мене пильнувати на цій дорозі, якою ходжу, і дасть мені хліба їсти та одежу вдягнутись,
GEN|28|21|і я з миром вернуся до дому батька свого, то Господь буде мені Богом,
GEN|28|22|і цей камінь, що я поставив за пам'ятника, буде домом Божим. І зо всього, що даси Ти мені, я, щодо десятини, дам десятину Тобі!
GEN|29|1|І зібрався Яків, і пішов до краю синів Кедему.
GEN|29|2|І побачив, аж ось криниця в полі, і ото там три отарі лежали біля неї, бо з тієї криниці напувають стада. А на отворі криниці лежав великий камінь.
GEN|29|3|І збирались туди всі стада, і скочували каменя з отвору криниці, і напоювали отару, і привалювали каменя на отвір криниці знов на його місце.
GEN|29|4|І сказав до пастухів Яків: Браття мої, звідкіля ви? А ті відказали: Ми з Харану.
GEN|29|5|І сказав їм: Чи ви знаєте Лавана, сина Нахорового? І відказали: Знаємо.
GEN|29|6|І сказав їм: Чи гаразд із ним? І відказали: Гаразд. А ось Рахіль, дочка його, приходить з отарою.
GEN|29|7|І сказав: Тож іще багато дня, не час зганяти худобу. Напійте отару, та йдіть пасіть.
GEN|29|8|А вони відказали: Не можемо, аж поки не будуть зігнані всі стада, і не відкотять каменя з отвору криниці, тоді понапуваємо отару.
GEN|29|9|Іще він говорив із ними, аж ось приходить Рахіль з отарою батька свого, бо була вона пастушка.
GEN|29|10|І сталося, коли Яків побачив Рахіль, дочку Лавана, брата своєї матері, то підійшов Яків і відкотив каменя з отвору криниці, і напоїв отару Лавана, брата матері своєї.
GEN|29|11|І поцілував Яків Рахіль, і підніс свій голос, і заплакав...
GEN|29|12|І Яків оповів Рахілі, що він брат батька її, і що він син Ревеки. А та побігла, і розповіла батькові своєму...
GEN|29|13|І сталося, коли Лаван почув вістку про Якова, сина сестри своєї, то побіг йому назустріч, і обняв його, і поцілував його, і привів його до свого дому. А він розповів Лаванові про всі ті пригоди.
GEN|29|14|І промовив до нього Лаван: Поправді, ти кість моя й тіло моє! І сидів він із ним місяць часу.
GEN|29|15|І сказав Лаван до Якова: Чи тому, що ти брат мій, то ти будеш служити мені даремно? Скажи ж мені, яка плата тобі?
GEN|29|16|А в Лавана було дві дочки: ім'я старшій Лія, а ім'я молодшій Рахіль.
GEN|29|17|Очі ж Ліїні були хворі, а Рахіль була гарного стану та вродливого вигляду.
GEN|29|18|І покохав Яків Рахіль, та й сказав: Я буду сім літ служити тобі за Рахіль, молодшу дочку твою.
GEN|29|19|І промовив Лаван: Краще мені віддати її тобі, аніж віддати мені її іншому чоловікові. Сиди ж зо мною!
GEN|29|20|І служив Яків за Рахіль сім літ, а вони через любов його до неї були в його очах, як кілька днів.
GEN|29|21|І сказав Яків Лаванові: Дай мені жінку мою, бо виповнилися мої дні, і нехай я до неї ввійду!
GEN|29|22|І зібрав Лаван усіх людей тієї місцевости, і справив гостину.
GEN|29|23|І сталося ввечері, і взяв він дочку свою Лію, і до нього впровадив її. І Яків із нею зійшовся.
GEN|29|24|А Лаван дав їй Зілпу, невільницю свою, дав Лії, дочці своїй, за невільницю.
GEN|29|25|А вранці виявилося, що то була Лія! І промовив Яків до Лавана: Що це ти вчинив мені? Хіба не за Рахіль працював я в тебе? Нащо ж обманив ти мене?
GEN|29|26|А Лаван відказав: У нашій місцевості не робиться так, щоб віддавати молодшу перед старшою.
GEN|29|27|Виповни тиждень для цієї, і буде дана тобі також та, за працю, що будеш працювати в мене ще сім літ других.
GEN|29|28|І зробив Яків так, і виповнив тиждень для цієї. І він дав йому Рахіль, дочку свою, дав йому за жінку.
GEN|29|29|І дав Лаван Рахілі, дочці своїй, Білгу, невільницю свою, дав їй за невільницю.
GEN|29|30|І прийшов він також до Рахілі, і покохав також Рахіль, більше, як Лію. І працював у нього ще сім літ других.
GEN|29|31|І побачив Господь, що зненавиджена Лія, і відкрив її утробу, а Рахіль була неплідна.
GEN|29|32|І завагітніла Лія, і сина породила, і назвала ім'я йому: Рувим, бо сказала була: Господь споглянув на недолю мою, бо тепер покохає мене чоловік мій!
GEN|29|33|І завагітніла вона ще, і сина породила, і сказала: Господь почув, що я зненавиджена, і дав мені також цього. І назвала ймення йому: Симеон.
GEN|29|34|І завагітніла вона ще, і сина породила, і сказала: Тепер оцим разом буде до мене прилучений мій чоловік, бо я трьох синів породила йому. Тому й назвала ім'я йому: Левій.
GEN|29|35|І завагітніла вона ще, і сина породила, і сказала: Тим разом я буду хвалити Господа! Тому назвала ім'я йому: Юда. Та й перестала роджати.
GEN|30|1|І побачила Рахіль, що вона не вродила Якову. І заздрила Рахіль сестрі своїй, і сказала до Якова: Дай мені синів! А коли ні, то я вмираю!
GEN|30|2|І запалився гнів Яковів на Рахіль, і він сказав: Чи я замість Бога, що затримав від тебе плід утроби?
GEN|30|3|І сказала вона: Ось невільниця моя Білга. Прийди до неї, і нехай вона вродить на коліна мої, і я також буду мати від неї дітей.
GEN|30|4|І вона дала йому Білгу, невільницю свою, за жінку. І ввійшов до неї Яків.
GEN|30|5|І завагітніла Білга, і вродила Якову сина.
GEN|30|6|І сказала Рахіль: Розсудив Бог мене, а також вислухав голос мій, і дав мені сина. Тому назвала ймення йому: Дан.
GEN|30|7|І завагітніла вона ще, і вродила Білга, невільниця Рахілина, другого сина Якову.
GEN|30|8|І сказала Рахіль: Великою боротьбою боролась я з сестрою своєю, і перемогла. І назвала ймення йому: Нефталим.
GEN|30|9|І побачила Лія, що вона перестала родити, і взяла Зілпу, свою невільницю, і дала її Якову за жінку.
GEN|30|10|І вродила Зілпа, невільниця Ліїна, Якову сина.
GEN|30|11|І сказала Лія: Прийшло щастя, і назвала ймення йому Ґад.
GEN|30|12|І вродила Зілпа, невільниця Ліїна, другого сина Якову.
GEN|30|13|І промовила Лія: То на блаженство моє, бо будуть уважати мене за жінку блаженну. І назвала ймення йому: Асир.
GEN|30|14|І пішов Рувим за тих днів, коли жато пшеницю, і знайшов на полі мандрагорові яблучка, і приніс їх до Лії, матері своєї. І сказала Рахіль до Лії: Дай мені з мандрагорових яблучок сина твого!
GEN|30|15|А та відказала їй: Чи мало тобі, що забрала мого чоловіка? І забереш також мандрагорові яблучка сина мого? І сказала Рахіль: Тому то він ляже з тобою цієї ночі за мандрагорові яблучка сина твого!
GEN|30|16|І прийшов Яків з поля ввечері, а Лія вийшла назустріч і сказала: Увійдеш до мене, бо справді найняла я тебе за мандрагорові яблучка сина мого. І лежав він із нею ночі тієї.
GEN|30|17|І вислухав Бог Лію, і завагітніла вона, і вродила Якову п'ятого сина.
GEN|30|18|І промовила Лія: Дав Бог заплату мені, що дала я невільницю свою своєму чоловікові. І назвала ймення йому: Іссахар.
GEN|30|19|І завагітніла Лія ще, і вродила Якову шостого сина.
GEN|30|20|І промовила Лія: Обдарував мене Бог добрим подарунком, цим разом замешкає в мене мій чоловік, бо я породила йому шестеро синів. І назвала ймення йому: Завулон.
GEN|30|21|А потому вродила дочку, і назвала ймення їй: Діна.
GEN|30|22|І згадав Бог про Рахіль, і вислухав її Бог, і відчинив їй утробу.
GEN|30|23|І завагітніла вона, і сина вродила, і сказала: Бог забрав мою ганьбу!
GEN|30|24|І назвала ймення йому: Йосип, кажучи: Додасть Господь мені іншого сина!
GEN|30|25|І сталося, коли Рахіль породила Йосипа, то сказав Яків до Лавана: Відпусти мене, і нехай я піду до свого місця й до Краю свого.
GEN|30|26|Дай же жінок моїх і дітей моїх, що служив тобі за них, і нехай я піду, бо ти знаєш службу мою, яку я служив був тобі.
GEN|30|27|І промовив до нього Лаван: Коли я знайшов милість в очах твоїх, побудь з нами, бо я зрозумів, що поблагословив мене Господь через тебе.
GEN|30|28|І далі казав: Признач собі заплату від мене, і я дам.
GEN|30|29|А той відказав: Ти знаєш, як я служив тобі, і якою стала худоба твоя зо мною.
GEN|30|30|Бо те мале, що було в тебе до мене, розмножилося на велике, і Господь поблагословив тебе, відколи нога моя в тебе. А тепер, коли ж я буду працювати для власного дому?
GEN|30|31|І сказав Лаван: Що ж я тобі дам? А Яків промовив: Не давай мені нічого. Коли зробиш мені оцю річ, то вернуся, буду пасти отару твою, буду пильнувати.
GEN|30|32|Я сьогодні перейду через усю отару твою, щоб вилучити звідти кожну овечку крапчасту й переполасу, і кожну овечку чорну з-поміж овець, і переполасе й крапчасте з-поміж кіз, і це буде заплата мені.
GEN|30|33|І справедливість моя посвідчить за мене в завтрішнім дні, коли прийдеш глянути на заплату мою від тебе. Усе, що воно не крапчасте й не переполасе з-поміж кіз і не чорне з-поміж овець, крадене воно в мене.
GEN|30|34|А Лаван відказав: Так, нехай буде за словом твоїм!
GEN|30|35|І того дня вилучив він козлів пасастих і покрапованих, і всі кози крапчасті й переполасі, усе, що біле було в ньому, і все чорне серед овець, і дав до рук своїх синів.
GEN|30|36|І визначив дорогу триденну поміж собою й поміж Яковом. А Яків пас позосталу Лаванову отару.
GEN|30|37|І взяв собі Яків сирого кия тополевого, і мігдалового, і каштанового, і налупив з них білих лушпин, відкриваючи білість, що на киях була.
GEN|30|38|І поставив кийки, що їх облупив, перед отарою при жолобах при коритах води, куди отара приходить пити. І вони злучувалися, як приходили пити.
GEN|30|39|І злучувалася отара при киях, і котилася овечками та козами пасастими, крапчастими й переполасими.
GEN|30|40|І відділяв Яків тих овечок, і ставив отару обличчям до пасастого й до всього чорного серед отари Лавана. І клав свої стада окремо, і не клав їх до отари Лаванової.
GEN|30|41|І бувало, що кожного разу, коли злучувалася отара міцна, то Яків клав при жолобах киї перед очі отари, щоб вона злучувалася при тих киях.
GEN|30|42|А як отара слаба була, то не клав. І ставалось, що слабе припадало Лаванові, а міцніше Якову.
GEN|30|43|І дуже-дуже зможнів той чоловік. І було в нього багато отар, і невільниці, і раби, і верблюди, і осли.
GEN|31|1|І почув був Яків слова Лаванових синів, що казали: Яків забрав усе, що було в нашого батька. І з того, що було в батька нашого, зробив собі всю оцю честь...
GEN|31|2|І побачив Яків Лаванове обличчя, а ото він тепер інший до нього, як був учора, позавчора.
GEN|31|3|І промовив Господь до Якова: Вернися до краю батьків своїх, і до місця твого народження. А Я буду з тобою.
GEN|31|4|І послав Яків, і покликав Рахіль і Лію на поле до отари своєї,
GEN|31|5|та й промовив до них: Я бачив обличчя вашого батька, що він тепер інший до мене, як був учора й позавчора. Та Бог батька мого був зо мною.
GEN|31|6|А ви знаєте, що всією силою своєю я служив вашому батькові.
GEN|31|7|І батько ваш сміявся з мене, і десять раз міняв заплату мені, але Бог не дав йому чинити зо мною зле.
GEN|31|8|Коли він говорив був отак: Крапчасте буде заплата твоя, то й котяться всі овечки та кози крапчасті. А коли скаже так: Пасасте буде заплата твоя, то й котяться всі овечки та кози пасасті.
GEN|31|9|І відняв Бог худобу вашого батька, та й дав мені.
GEN|31|10|І сталося в час, коли отара злучувалася, звів був я очі свої та й побачив у сні: аж ось козли, що спинались на овечок та на кіз, були пасасті, крапчасті й рябі.
GEN|31|11|І сказав мені Ангол у сні: Якове! А я відказав: Ось я!
GEN|31|12|Він промовив: Зведи свої очі й побач: усі козли, що спинаються на овечок та на кіз, пасасті, крапчасті й рябі, бо Я бачив усе, що Лаван виробляє тобі.
GEN|31|13|Я Бог Бет-Елу, що ти намастив був там пам'ятника, і Мені склав там обітницю. Тепер уставай, вийди з цієї землі, і вертайся до землі твого народження.
GEN|31|14|І відповіла Рахіль та Лія, та й сказали йому: Чи ми маємо частку та спадщину в домі нашого батька?
GEN|31|15|Таж він нас полічив за чужинців, бо продав нас, і справді пожер наше срібло.
GEN|31|16|Бож усе багатство, що Бог вирвав від нашого батька, воно наше та наших синів. А тепер зроби все, що Бог наказав був тобі.
GEN|31|17|І встав Яків, і посадив синів своїх і жінок своїх на верблюди.
GEN|31|18|І він забрав усю худобу свою, і все майно своє, що набув, здобуту худобу свою, що набув у Падані арамейськім, щоб прийти до Ісака, батька свого, до землі ханаанської.
GEN|31|19|А Лаван пішов стригти отару свою, а Рахіль покрала домових божків, яких батько мав.
GEN|31|20|І Яків обманив Лавана арамейського, бо не сказав йому, що втікає.
GEN|31|21|І втік він, і все, що його. І встав, і перейшов річку, і прямував до Ґілеядської гори.
GEN|31|22|А третього дня розказано Лаванові, що Яків утік.
GEN|31|23|І взяв він з собою братів своїх, і гнався за ним дорогою семи день, та й догнав його на горі Ґілеядській.
GEN|31|24|І прийшов Бог до Лавана арамеянина в нічнім сні, та й до нього сказав: Стережися, щоб ти не говорив з Яковом ані доброго, ані злого.
GEN|31|25|І догнав Лаван Якова. А Яків поставив намета свого на горі, і Лаван поставив з братами своїми на горі Ґілеядській.
GEN|31|26|І промовив Лаван до Якова: Що ти зробив? Ти обманив мене, і забрав моїх дочок, немов бранок меча!
GEN|31|27|Чого втік ти таємно, і обікрав мене, і не сказав мені? А я був би відіслав тебе з радістю, із співами, з бубном, і з гуслами.
GEN|31|28|І ти не дозволив мені навіть поцілувати онуків моїх і дочок моїх. Тож ти нерозумно вчинив!
GEN|31|29|Я маю в руці своїй силу, щоб учинити з вами зле. Але Бог вашого батька вчора вночі сказав був до мене, говорячи: Стережися, щоб ти не говорив з Яковом ані доброго, ані злого.
GEN|31|30|А тепер справді підеш, бо ти сильно затужив за домом батька свого. Але нащо ти покрав моїх богів?
GEN|31|31|А Яків відповів і сказав до Лавана: Тому, що боявся, бо я думав: Аби но він не забрав від мене своїх дочок!
GEN|31|32|При кому ж ти знайдеш своїх богів, не буде він жити. Перед нашими братами пізнай собі, що твого в мене, і візьми собі. А Яків не знав, що Рахіль їх покрала.
GEN|31|33|І ввійшов Лаван до намету Якового, і до намету Ліїного, і до намету обох невільниць, та нічого не знайшов. І вийшов він із намету Ліїного і ввійшов до намету Рахілиного.
GEN|31|34|А Рахіль узяла божки, і вложила їх до сідла верблюда, та й сіла на них. І обмацав Лаван усього намета, і нічого не знайшов.
GEN|31|35|А вона сказала до батька свого: Нехай не палає гнів в очах батька мого, бо я не можу встати перед обличчям твоїм, бо в мене тепер звичайне жіноче. І перешукав він, та божків не знайшов.
GEN|31|36|І запалав Яків гнівом, і сварився з Лаваном. І відповів Яків, і сказав до Лавана: Яка провина моя, який мій гріх, що ти гнався за мною,
GEN|31|37|що ти обмацав усі мої речі? Що ти знайшов зо всіх речей свого дому, положи тут перед моїми братами і братами своїми, і нехай вони розсудять поміж нами двома.
GEN|31|38|Я вже двадцять літ із тобою. Вівці твої та кози твої не мертвили свого плоду, а баранів отари твоєї я не їв.
GEN|31|39|Розшарпаного диким звірем я не приносив до тебе, я сам ніс ту шкоду. Від мене домагався ти того, що було вкрадене вдень, і що було вкрадене вночі.
GEN|31|40|Бувало, що вдень з'їдала мене спекота, а вночі паморозь, а мій сон мандрував від моїх очей.
GEN|31|41|Таке мені двадцять літ у твоїм домі... Служив я тобі чотирнадцять літ за двох дочок твоїх, і шість літ за отару твою, а ти десять раз зміняв мені свою заплату!
GEN|31|42|Коли б не був при мені Бог батька мого, Бог Авраамів, і не Той, Кого боїться Ісак, то тепер ти відіслав би мене впорожні!... Біду мою й труд рук моїх Бог бачив, і виказав це вчора вночі.
GEN|31|43|І відповів Лаван і сказав до Якова: Дочки дочки мої, а діти мої діти, а отара моя отара, і все, що ти бачиш то моє. А дочкам моїм, що зроблю їм сьогодні, або їхнім дітям, що вони породили їх?
GEN|31|44|А тепер ходи, я й ти вчинімо умову, і оце буде свідком поміж мною й поміж тобою.
GEN|31|45|І взяв Яків каменя, і поставив його за пам'ятника.
GEN|31|46|І сказав Яків браттям своїм: Назбирайте каміння. І назбирали каміння вони, та й зробили могилу, і їли там на тій могилі.
GEN|31|47|І назвав її Лаван: Еґар-Сагадута, а Яків її назвав: Ґал-Ед.
GEN|31|48|І промовив Лаван: Ця могила свідок між мною й між тобою сьогодні, тому то й названо ймення її: Ґал-Ед
GEN|31|49|і Міцпа, бо сказав: Нехай дивиться Господь між мною й між тобою, коли ми розійдемося один від одного.
GEN|31|50|Коли ти будеш кривдити дочок моїх, і коли візьмеш за жінок понад дочок моїх, то не людина з нами, а дивися Бог свідок між мною й між тобою!
GEN|31|51|А Яків сказав до Лавана: Ось ця могила, й ось той пам'ятник, якого поставив я між собою й між тобою.
GEN|31|52|Свідок ця могила, і свідок цей пам'ятник, що я не перейду цієї могили до тебе, і ти не перейдеш до мене цієї могили та цього пам'ятника на зле.
GEN|31|53|Розсудить між нами Бог Авраамів і Бог Нахорів, Бог їхнього батька. І Яків присягнув Тим, Кого боїться його батько Ісак.
GEN|31|54|І приніс Яків жертву на горі, і покликав братів своїх їсти хліб. І вони їли хліб і ночували на горі.
GEN|31|55|(32-1) І встав Лаван рано вранці, і поцілував онуків своїх, і дочок своїх, і поблагословив їх. І пішов, та й вернувся Лаван до місця свого.
GEN|32|1|(32-2) А Яків пішов на дорогу свою. І спіткали його Божі Анголи.
GEN|32|2|(32-3) І Яків сказав, коли їх побачив: Це Божий табір! І він назвав ім'я тому місцю: Маханаїм.
GEN|32|3|(32-4) І послав Яків послів перед собою до Ісава, брата свого, до землі Сеїр, до краю едомського.
GEN|32|4|(32-5) І наказав їм, говорячи: Скажіть так моєму панові Ісавові: Так сказав раб твій Яків: Я мешкав з Лаваном, і задержався аж дотепер.
GEN|32|5|(32-6) І маю я вола та осла, і отару, і раба, і невільницю. І я послав розказати панові моєму, щоб знайти милість в очах твоїх.
GEN|32|6|(32-7) І вернулися посли до Якова, та й сказали: Ми прийшли були до брата твого до Ісава, а він також іде назустріч тобі, і чотири сотні людей з ним.
GEN|32|7|(32-8) І Яків сильно злякався, і був затурбований. І він поділив народ, що був з ним, і дрібну та велику худобу, і верблюди на два табори.
GEN|32|8|(32-9) І сказав: Коли прийде Ісав до табору одного, і розіб'є його, то вціліє позосталий табір.
GEN|32|9|(32-10) І Яків промовив: Боже батька мого Авраама, і Боже батька мого Ісака, Господи, що сказав Ти мені: Вернися до Краю свого, і до місця свого народження, і Я зроблю тобі добре.
GEN|32|10|(32-11) Я не вартий усіх отих милостей, і всієї вірности, яку Ти чинив був Своєму рабові, бо з самою своєю палицею перейшов я був цей Йордан, а тепер я стався на два табори.
GEN|32|11|(32-12) Збережи ж мене від руки мого брата, від руки Ісава, бо боюсь я його, щоб він не прийшов та не побив мене і матері з дітьми.
GEN|32|12|(32-13) А Ти ж був сказав: Учинити добро учиню я з тобою добро; а нащадки твої покладу, як той морський пісок, що його не злічити через безліч.
GEN|32|13|(32-14) І він переночував там тієї ночі, і взяв із того, що під руку прийшло, дар для Ісава, брата свого:
GEN|32|14|(32-15) кіз двісті, і козлів двадцятеро, овець двісті, і баранів двадцятеро,
GEN|32|15|(32-16) верблюдиць дійних та їх жереб'ят тридцятеро, корів сорок, а биків десятеро, ослиць двадцятеро, а ослят десятеро.
GEN|32|16|(32-17) І дав до рук рабів своїх кожне стадо окремо. І сказав він до рабів своїх: Ідіть передо мною, і позоставте відстань поміж стадом і стадом.
GEN|32|17|(32-18) І він наказав першому, кажучи: Коли спіткає тебе Ісав, брат мій, і запитає тебе так: Чий ти, і куди ти йдеш, і чиє те, що перед тобою?
GEN|32|18|(32-19) то скажеш: Раба твого Якова це подарунок, посланий панові моєму Ісавові. А ото й він сам за нами.
GEN|32|19|(32-20) І наказав він і другому, і третьому, також усім, що йшли за стадами, говорячи: Таким словом будете говорити до Ісава, коли ви знайдете його,
GEN|32|20|(32-21) і скажете: Ось і раб твій Яків за нами, бо він сказав: Нехай я вблагаю його оцим дарунком, що йде передо мною, а потім побачу обличчя його, може він підійме обличчя моє.
GEN|32|21|(32-22) І йшов подарунок перед ним, а він ночував тієї ночі в таборі.
GEN|32|22|(32-23) І встав він тієї ночі, і взяв обидві жінки свої, і обидві невільниці свої та одинадцятеро дітей своїх, і перейшов брід Яббок.
GEN|32|23|(32-24) І він узяв їх, і перепровадив через потік, і перепровадив те, що в нього було.
GEN|32|24|(32-25) І зостався Яків сам. І боровся з ним якийсь Муж, аж поки не зійшла досвітня зоря.
GEN|32|25|(32-26) І Він побачив, що не подужає його, і доторкнувся до суглобу стегна його. І звихнувся суглоб стегна Якова, як він боровся з Ним.
GEN|32|26|(32-27) І промовив: Пусти Мене, бо зійшла досвітня зоря. А той відказав: Не пущу Тебе, коли не поблагословиш мене.
GEN|32|27|(32-28) І промовив до нього: Як твоє ймення? Той відказав: Яків.
GEN|32|28|(32-29) І сказав: Не Яків буде називатися вже ймення твоє, але Ізраїль, бо ти боровся з Богом та з людьми, і подужав.
GEN|32|29|(32-30) І запитав Яків і сказав: Скажи ж Ім'я Своє. А Той відказав: Пощо питаєш про Ймення Моє? І Він поблагословив його там.
GEN|32|30|(32-31) І назвав Яків ім'я того місця: Пенуїл, бо бачив був Бога лицем у лице, та збереглася душа моя.
GEN|32|31|(32-32) І засвітило йому сонце, коли він перейшов Пенуїл. І він кульгав на своє стегно.
GEN|32|32|(32-33) Тому не їдять Ізраїлеві сини жили стегна, що на суглобі стегна, аж до сьогодні, бо Він доторкнувся був до стегна Якового, жили стегна.
GEN|33|1|І звів Яків очі свої, та й побачив, аж ось іде Ісав, а з ним чотири сотні людей. І він поділив своїх дітей на Лію, і на Рахіль, і на обох невільниць своїх.
GEN|33|2|І поставив він тих невільниць і дітей їх напереді, а Лію й дітей її передостанніми, а Рахіль та Йосипа останніми.
GEN|33|3|А сам пішов перед ними, і вклонився до землі сім раз, аж поки підійшов до брата свого.
GEN|33|4|І побіг Ісав назустріч йому, і обняв його, і впав на шию йому, і цілував його. І вони заплакали.
GEN|33|5|І звів свої очі Ісав, і побачив жінок та дітей. І сказав: Хто то такі? А той відказав: Діти, якими обдарував Бог твого раба.
GEN|33|6|І підійшли сюди невільниці, і їхні діти, та й вклонилися.
GEN|33|7|І підійшла також Лія та діти її, і вклонилися, а потім підійшов Йосип і Рахіль, та й вклонилися.
GEN|33|8|І сказав Ісав: А що це за цілий табір той, що я спіткав? А той відказав: Щоб знайти милість в очах мого пана.
GEN|33|9|А Ісав сказав: Я маю багато, мій брате, твоє нехай буде тобі.
GEN|33|10|А Яків сказав: Ні ж бо! Коли я знайшов милість в очах твоїх, то візьми дарунка мого з моєї руки. Бож я побачив обличчя твоє, ніби побачив Боже лице, і ти собі уподобав мене.
GEN|33|11|Візьми ж благословення моє, що припроваджене тобі, бо Бог був милостивий до мене, та й маю я все. І благав він його, і той узяв.
GEN|33|12|І промовив Ісав: Рушаймо й ходім, а я піду обік тебе.
GEN|33|13|А той відказав: Пан мій знає, що діти молоді, а дрібна та велика худоба в мене дійні. Коли погнати їх один день, то вигине вся отара.
GEN|33|14|Нехай же піде пан мій перед очима свого раба, а я піду поволі за ногою скотини, що передо мною, і за ногою дітей, аж поки не прийду до пана свого до Сеїру.
GEN|33|15|І промовив Ісав: Позоставлю ж з тобою трохи з людей, що зо мною. А той відказав: Пощо знаходжу я таку милість в очах свого пана?.
GEN|33|16|І вернувся того дня Ісав на дорогу свою до Сеїру.
GEN|33|17|А Яків подався до Суккоту, і збудував собі хату, а для худоби своєї поробив курені, тому назвав ім'я тому місцю: Суккот.
GEN|33|18|І Яків, коли він прийшов із Падану арамейського, прибув спокійно до міста Сихем у Краї ханаанському, і розтаборився перед містом.
GEN|33|19|І купив він кусок поля, де розклав намета свого, з руки синів Гамора, батька Сихема, за сто срібняків.
GEN|33|20|І поставив там жертівника, і назвав його: Ел-Елогей-Ізраїль.
GEN|34|1|І вийшла була Діна, дочка Лії, яка вродила її Якову, щоб подивитися на дочок того краю.
GEN|34|2|І побачив її Сихем, син Гамора хівеянина, начальника того краю, і взяв її, і лежав із нею, і збезчестив її.
GEN|34|3|І пригорнулася душа його до Діни, дочки Якової, і покохав він дівчину, і говорив до серця дівочого.
GEN|34|4|І сказав Сихем до Гамора, батька свого, говорячи: Візьми те дівча за жінку для мене!
GEN|34|5|А Яків почув, що той збезчестив Діну, дочку його, а сини його були з худобою його на полі. І мовчав Яків, аж поки прибули вони.
GEN|34|6|І вийшов Гамор, Сихемів батько, до Якова, щоб поговорити з ним.
GEN|34|7|І прийшли сини Яковові з поля, коли почули, і засмутились ці люди, і сильно запалав їхній гнів, бо той ганьбу зробив в Ізраїлі тим, що лежав із дочкою Якова, а так не робиться.
GEN|34|8|А Гамор говорив з ними, кажучи: Син мій Сихем, запрагла душа його вашої дочки. Дайте ж її йому за жінку!
GEN|34|9|І посвоячтеся з нами, дайте нам ваші дочки, а наші дочки візьміть собі.
GEN|34|10|І осядьтеся з нами, а цей край буде перед вами. Сидіть і перемандруйте його, і набувайте на власність у нім.
GEN|34|11|І промовив Сихем до батька її та до братів її: Нехай я знайду милість у ваших очах, і що ви скажете мені я дам.
GEN|34|12|Сильно побільшіть на мене віно та дарунок, а я дам, як мені скажете, та тільки дайте мені дівчину за жінку!
GEN|34|13|І відповіли сини Якова Сихемові та Гаморові, батькові його, підступом, сказали, бо він збезчестив Діну, сестру їх.
GEN|34|14|І сказали до них: Ми не можемо зробити тієї речі, видати сестру нашу чоловікові, що має крайню плоть, бо то ганьба для нас.
GEN|34|15|Ми тільки за те прихилимось до вас, коли ви станете, як ми, щоб у вас був обрізаний кожний чоловічої статі.
GEN|34|16|І дамо вам своїх дочок, а ваших дочок візьмемо собі, й осядемось із вами, і станемо одним народом.
GEN|34|17|А коли ви не послухаєте нас, щоб обрізатися, то ми візьмемо свої дочки, та й підемо.
GEN|34|18|І їхні слова були добрі в очах Гамора та в очах Сихема, сина Гаморового.
GEN|34|19|І не загаявся юнак той учинити ту річ, бо полюбив дочку Якова. А він був найповажніший у всім домі батька свого.
GEN|34|20|І прибув Гамор та Сихем, син його, до брами міста, і промовили до людей свого міста, говорячи:
GEN|34|21|Ці люди вони приязні до нас, і нехай осядуть у краю, і нехай перемандрують його, а цей край ось розлогий перед ними. Дочок їхніх візьмімо собі за жінок, а наших дочок даймо їм.
GEN|34|22|Тільки за це прихиляться до нас ці люди, щоб сидіти з нами, і щоб стати одним народом, коли в нас буде обрізаний кожен чоловічої статі, як і вони обрізані.
GEN|34|23|Отара їхня, і майно їхнє, і вся їхня худоба хіба не наші вони? Тільки прихилімося до них, і нехай вони осядуть із нами.
GEN|34|24|І послухали Гамора та Сихема, сина його, усі, хто виходив з брами його міста. І були обрізані всі чоловічої статі, усі, хто виходив з брами міста його.
GEN|34|25|І сталося третього дня, коли вони хворі були, то два сини Яковові, Симеон і Левій, брати Дінині, взяли кожен меча свого, і безпечно напали на місто, і повбивали всіх чоловіків.
GEN|34|26|Також Гамора й Сихема, сина його, забили мечем, і забрали Діну з дому Сихемового, та й вийшли.
GEN|34|27|Сини Якова напали на трупи, і пограбували місто за те, що вони збезчестили їхню сестру.
GEN|34|28|Забрали дрібну й велику худобу їх, і осли їх, і що було в місці, і що на полі,
GEN|34|29|і ввесь маєток їхній, і всіх їхніх дітей, і їхніх жінок забрали в неволю, і пограбували все, що де в домі було.
GEN|34|30|І сказав Яків до Симеона й до Левія: Ви зробили мене нещасливим, бо зробили мене зненавидженим у мешканців цього краю, у ханаанеянина й периззеянина. Ми люди нечисленні, а вони зберуться на мене, та й поб'ють мене, і буду знищений я та мій дім.
GEN|34|31|А вони відказали: Чи він мав би зробити нашу сестру блудницею?
GEN|35|1|І сказав Бог до Якова: Уставай, вийди до Бет-Елу, і там осядься, і зроби там жертівника Богові, що явився тобі, як ти втікав був перед Ісавом, братом своїм.
GEN|35|2|І сказав Яків до дому свого, до всіх, хто був із ним: Усуньте чужинних богів, які є серед вас, і очистьтеся, і змініть свою одіж.
GEN|35|3|І встаньмо, і підім до Бет-Елу, і зроблю я там жертівника Богові, що відповів мені в день мого утиску, і був зо мною в дорозі, якою ходив я.
GEN|35|4|І вони віддали Якову всіх чужинних богів, що були в їх руках, і сережки, що в їхніх ушах, а Яків сховав їх під дубом, що перед Сихемом.
GEN|35|5|І вирушили вони. І великий жах обгорнув ті міста, що навколо них, і вони не гналися за синами Якова.
GEN|35|6|І прибув Яків до Лузу, що в землі ханаанській, цебто до Бет-Елу, він і ввесь народ, що був з ним.
GEN|35|7|І збудував він там жертівника, та й назвав те місце: Ел Бет-Ел, бо там явився йому Бог, коли він утікав перед своїм братом.
GEN|35|8|І вмерла Девора, мамка Ревеки, і була похована нижче Бет-Елу під дубом, а він назвав ім'я йому: Аллон-Бахут.
GEN|35|9|І ще явився Бог до Якова, коли він прийшов був із Падану арамейського, і поблагословив його.
GEN|35|10|І сказав йому Бог: Ім'я твоє Яків. Не буде вже кликатися ім'я твоє Яків, але Ізраїль буде ім'я твоє. І назвав ім'я йому: Ізраїль.
GEN|35|11|І сказав йому Бог: Я Бог Всемогутній! Плодися й розмножуйся, народ і громада народів буде з тебе, і царі вийдуть із стегон твоїх.
GEN|35|12|А той Край, що я дав його Авраамові та Ісакові, дам його тобі, і нащадку твоєму по тобі дам Я той Край.
GEN|35|13|І вознісся Бог з-понад нього в місці, де з ним говорив.
GEN|35|14|І поставив Яків пам'ятника на тому місці, де Він говорив з ним, пам'ятника кам'яного, і вилив на нього винне лиття, і полив його оливою.
GEN|35|15|І назвав Яків ім'я місцю, що там говорив із ним Бог: Бет-Ел.
GEN|35|16|І він рушив із Бет-Елу. І була ще ківра землі до Ефрати, а Рахіль породила, і були важкі її пологи.
GEN|35|17|І сталося, коли важкі були її пологи, то сказала їй баба-сповитуха: Не бійся, бо й це тобі син.
GEN|35|18|І сталося, коли виходила душа її, бо вмирала вона, то назвала ім'я йому: Бен-Оні, а його батько назвав його: Веніямин.
GEN|35|19|І вмерла Рахіль, і була похована на дорозі до Ефрати, це є Віфлеєм.
GEN|35|20|І поставив Яків пам'ятника на гробі її, це надгробний пам'ятник Рахілі аж до сьогодні.
GEN|35|21|І рушив Ізраїль, і розтягнув намета свого далі до Міґдал-Едеру.
GEN|35|22|І сталося, коли Ізраїль перебував у тім краї, то Рувим пішов і ліг із Білгою, наложницею батька свого. І почув Ізраїль, і було це злим йому. А в Якова було дванадцятеро синів.
GEN|35|23|Сини Ліїні: перворідний Якова Рувим, і Симеон, і Левій, і Юда, і Іссахар, і Завулон.
GEN|35|24|Сини Рахілині: Йосип і Веніямин.
GEN|35|25|А сини Білги, невільниці Рахілиної: Дан і Нефталим.
GEN|35|26|А сини Зілпи, невільниці Ліїної: Ґад і Асир. Оце сини Якова, що йому народжено в Падані арамейському.
GEN|35|27|І прибув Яків до Ісака, свого батька, до Мамре, до Кир'ят-Арби, цебто Хеврону, що там жив Авраам та Ісак.
GEN|35|28|І були Ісакові дні сто літ і вісімдесят літ.
GEN|35|29|І впокоївся Ісак та й помер, і прилучився до своєї рідні, старий та нажившись. І поховали його Ісав та Яків, сини його.
GEN|36|1|А оце нащадки Ісава, цебто Едома.
GEN|36|2|Ісав узяв жінок своїх з дочок ханаанських, Аду, дочку Елона хіттеянина, та Оголіваму, дочку Ани, дочку Ців'она хівеянина,
GEN|36|3|та Босмат, дочку Ізмаїлову, сестру Невайотову.
GEN|36|4|І породила Ада Ісавові Еліфаза, а Босмат породила Реуїла,
GEN|36|5|а Оголівама породила Суша, і Ялама, і Кораха. Оце сини Ісавові, що були йому народжені в ханаанській землі.
GEN|36|6|І взяв Ісав жінок своїх, і синів своїх, і дочок своїх, і всі душі дому свого, і худобу свою, і все стадо своє, і все своє майно, що набув у ханаанській землі, та й пішов до Краю від обличчя Якова, брата свого,
GEN|36|7|бо маєток їх був більший, щоб пробувати їм разом, і край їх часового замешкання не міг вмістити їх через їхню худобу.
GEN|36|8|І осівся Ісав на горі Сеїр, Ісав він Едом.
GEN|36|9|А оце нащадки Ісава, батька Едому на горі Сеїр.
GEN|36|10|Оце ймення синів Ісавових: Еліфаз, син Ади, жінки Ісавової, Реуїл, син Босмати, Ісавової жінки.
GEN|36|11|А сини Еліфазові були: Теман, Омар, Цефо, і Ґатам, і Кеназ.
GEN|36|12|А Тимна була наложниця Еліфаза, Ісавового сина, і породила вона Еліфазові Амалика. Оце сини Ади, Ісавової жінки.
GEN|36|13|А оце сини Реуїлові: Нагат і Зера, Шамма й Мізза. Оце сини Босмати, Ісавової жінки.
GEN|36|14|А оці були сини Оголівами, дочки Ани, дочки Ців'она, Ісавової жінки, і вродила вона Ісаву, Єуша, і Ялама, і Корея.
GEN|36|15|А оце провідники Ісавових синів. Сини Еліфаза, Ісавового перворідного: провідник Теман, провідник Омар, провідник Цефо, провідник Кеназ,
GEN|36|16|провідник Корей, провідник Ґатам, провідник Амалик. Оце провідники Еліфаза в краю Едома, оце сини Ади.
GEN|36|17|А оце сини Реуїла, Ісавового сина: провідник Нагат, провідник Зерах, провідник Шамма, провідник Мізза. Оце провідники Реуїлові в краю едомському, оце сини Босмати, Ісавової жінки.
GEN|36|18|А оце сини Оголівами, жінки Ісава: провідник Еуш, провідник Ялам, провідник Корей, оце провідники Оголівами, дочки Ани, Ісавової жінки.
GEN|36|19|Оце сини Ісава, цебто Едома, і оце їхні провідники.
GEN|36|20|Оце сини Сеїра, хореянина, мешканці цієї землі: Лотан і Шовал, і Ців'он, і Ана,
GEN|36|21|і Дішон, і Ецев, і Дішан, оце провідники хореянина, сини Сеїру, краю едомського.
GEN|36|22|А сини Лотана були: Хорі й Гемам, а Лотанова сестра Тимна.
GEN|36|23|А оце сини Шовалові: Алван і Манахат, і Евал, Шефо, і Онам.
GEN|36|24|А ото сини Ців'онові: і Айя, і Ана, той Ана, що знайшов був в пустині гарячі джерела, коли пас осли Ців'она, свого батька.
GEN|36|25|А оце діти Ани: Дішон, і Оголівама, дочка Ани.
GEN|36|26|А оце сини Дішонові: Хемдан, і Ешбан, і Ітран, і Керан.
GEN|36|27|Ото сини Ецера: Білган, і Зааван, і Акан.
GEN|36|28|Оце сини Дішана: Уц і Аран.
GEN|36|29|Оце провідники хореянина: провідник Лотан, провідник Шовал, провідник Ців'он, провідник Ана,
GEN|36|30|провідник Дішон, провідник Ецер, провідник Дішан, оце провідники хореянина за їхніми провідниками в краї Сеїр.
GEN|36|31|А оце царі, що царювали в краю Едома перед царюванням царя в синів Ізраїлевих.
GEN|36|32|І царював в Едомі Бела, син Беора, а ймення його міста Дінгава.
GEN|36|33|І вмер Бела, і зацарював замість нього Йовав, син Зераха з Боцри.
GEN|36|34|І вмер Йовав, і зацарював замість нього Хушам із землі теманіянина.
GEN|36|35|І вмер Хушам, і зацарював замість нього Гадад, син Бедада, що побив мідіян на полі Моава, а ймення його міста Авіт.
GEN|36|36|І вмер Гадад, і зацарював замість нього Самла з Машеку.
GEN|36|37|І вмер Самла, і зацарював замість нього Саул з Реховоту надрічного.
GEN|36|38|І вмер Саул, і зацарював замість нього Баал-Ханан, син Ахборів.
GEN|36|39|І вмер Баал-Ханан, син Ахборів, і зацарював замість нього Гадад, а ім'я його міста Пау, а ім'я його жінки Мегетав'іл, дочка Матреди, дочки Ме-Загава.
GEN|36|40|А оце імена провідників Ісавових за їхніми родами, за місцями їх, їхніми іменами: провідник Тимна, провідник Алва, провідник Етет,
GEN|36|41|провідник Оголівама, провідник Ела, провідник Пінон,
GEN|36|42|провідник Кеназ, провідник Теман, провідник Мівцар,
GEN|36|43|провідник Маґдіїл, провідник Ірам. Оце провідники Едома він же Ісав, батько Едому за їхніми оселями в краї їхнього володіння.
GEN|37|1|І осівся Яків у Краї мешкання батька свого, в Краї ханаанському.
GEN|37|2|Оце оповість про Якова. Йосип, віку сімнадцяти літ, пас, як юнак, отару з братами своїми, з синами Білги та з синами Зілпи, жінок батька свого. І Йосип доносив недобрі звістки про них до їхнього батька.
GEN|37|3|А Ізраїль любив Йосипа над усіх синів своїх, бо він був у нього сином старости. І він справив йому квітчасте вбрання.
GEN|37|4|І бачили його браття, що їх батько полюбив його над усіх братів його, і зненавиділи його, і не могли говорити з ним спокійно.
GEN|37|5|І снився був Йосипові сон, і він розповів своїм браттям, а вони ще збільшили ненависть до нього.
GEN|37|6|І сказав він до них: Послухайте но про той сон, що снився мені.
GEN|37|7|А ото ми в'яжемо снопи серед поля, і ось мій сніп зачав уставати, та й став. І ось оточують ваші снопи, та й вклоняються снопові моєму.
GEN|37|8|І сказали йому його браття: Чи справді ти будеш царювати над нами, чи теж справді ти будеш панувати над нами? І вони збільшили ненависть до нього через сни його та через слова його.
GEN|37|9|І снився йому ще сон інший, і він оповів його братам своїм, та й сказав: Оце снився мені ще сон, і ось сонце та місяць та одинадцять зір вклоняються мені.
GEN|37|10|І він розповів це батькові своєму та браттям своїм. І докорив йому батько його, та й промовив до нього: Що то за сон, що снився тобі? Чи справді прийдемо ми, я та мати твоя та брати твої, щоб уклонитися тобі до землі?
GEN|37|11|І заздрили йому брати його, а батько його запам'ятав ці слова.
GEN|37|12|І пішли брати його пасти отару свого батька в Сихем.
GEN|37|13|І сказав Ізраїль до Йосипа: Таж брати твої пасуть у Сихемі! Іди ж, і я пошлю тебе до них! А той відказав йому: Ось я!
GEN|37|14|І сказав він до нього: Піди но, побач стан братів твоїх і стан отари, та й дай мені відповідь. І він послав його з долини Хеврону, і той прибув до Сихему.
GEN|37|15|І знайшов його один чоловік, а він ось блукає по полю. І запитав його той чоловік, кажучи: Чого ти шукаєш?
GEN|37|16|А той відказав: Я шукаю братів своїх. Скажи ж мені, де вони випасають?
GEN|37|17|І сказав той чоловік: Вони пішли звідси, бо я чув, як казали вони: Ходімо до Дотаїну. І пішов Йосип за своїми братами, і знайшов їх у Дотаїні.
GEN|37|18|А вони побачили його здалека, і поки він наблизився до них, то змовлялися на нього, щоб убити його.
GEN|37|19|І сказали вони один одному: Ось іде той сновидець!
GEN|37|20|А тепер давайте вбиймо його, і вкиньмо його до однієї з ям, та й скажемо: Дикий звір з'їв його! І побачимо, що буде з його снами.
GEN|37|21|І почув це Рувим, і визволив його з руки їхньої, і сказав: Не губімо душі його!
GEN|37|22|І сказав до них Рувим: Не проливайте крови, киньте його до ями тієї, що в пустині, а руки не кладіть на нього, щоб визволити його з їхньої руки, щоб вернути його до батька його.
GEN|37|23|І сталося, коли прийшов Йосип до братів своїх, то вони стягнули з Йосипа вбрання його, вбрання квітчасте, що на ньому було.
GEN|37|24|І взяли його, та й кинули його до ями, а яма та порожня була, не було в ній води.
GEN|37|25|І сіли вони попоїсти хліба. І звели вони очі свої та й побачили, ось караван ізмаїлітів іде з Ґілеаду, а верблюди їхні несуть пахощі, і бальзам, і ладан, іде він спровадити це до Єгипту.
GEN|37|26|І сказав Юда до своїх братів: Яка користь, що вб'ємо нашого брата, і затаїмо його кров?
GEN|37|27|Давайте продамо його ізмаїльтянам, і рука наша нехай не буде на ньому, бо він брат нам, він наше тіло. І послухалися брати його.
GEN|37|28|І коли проходили мідіяніти, купці, то витягли й підняли Йосипа з ями. І продали Йосипа ізмаїльтянам за двадцять срібняків, а ті повели Йосипа до Єгипту.
GEN|37|29|А Рувим вернувся до ями, аж нема Йосипа в ямі! І розірвав він одежу свою...
GEN|37|30|І вернувся він до братів своїх, та й сказав: Немає хлопця! А я, куди я піду?
GEN|37|31|А вони взяли Йосипове вбрання, і зарізали козла, і вмочили вбрання в кров.
GEN|37|32|І послали вони квітчасте вбрання, і принесли до свого батька, та й сказали: Оце ми знайшли. Пізнай но, чи це вбрання твого сина воно, чи ні?
GEN|37|33|А він пізнав його та й сказав: Вбрання мого сина... Дикий звір його з'їв... Справді розшарпаний Йосип!
GEN|37|34|І роздер Яків одіж свою, і зодягнув веретище на стегна свої, і багато днів справляв жалобу по синові своєму...
GEN|37|35|І зачали всі сини його та всі дочки його потішати його. Але він не міг утішитися, та й сказав: У жалобі зійду я до сина мого до шеолу. І плакав за ним його батько.
GEN|37|36|І мідіяніти продали Йосипа до Єгипту, до Потіфара, царедворця фараонового, начальника царської сторожі.
GEN|38|1|Сталося того часу, і відійшов Юда від братів своїх, і розташувався аж до одного адулламітянина, а ймення йому Хіра.
GEN|38|2|І побачив там Юда дочку одного ханаанеянина, а ім'я йому Шуа, і взяв її, і з нею зійшовся.
GEN|38|3|І завагітніла вона, і породила сина, а він назвав ім'я йому: Ер.
GEN|38|4|І завагітніла вона ще, і породила сина, і назвала ім'я йому: Онан.
GEN|38|5|І ще знову, і породила сина, і назвала ім'я йому: Шела. А батько був у Кезиві, як вона породила його.
GEN|38|6|І взяв Юда жінку для Ера, свого перворідного, а ім'я їй: Тамара.
GEN|38|7|І був Ер, Юдин перворідний, злий в очах Господа, і Господь його вбив.
GEN|38|8|І сказав Юда до Онана: Увійди до жінки брата свого, і одружися з нею, і встанови насіння для брата свого.
GEN|38|9|А Онан знав, що не його буде насіння те. І сталося, коли він сходився з жінкою брата свого, то марнував насіння на землю, аби не дати його своєму братові.
GEN|38|10|І було зле в очах Господа те, що він чинив, і вбив Він також його.
GEN|38|11|І сказав Юда до Тамари, невістки своєї: Сиди вдовою в домі батька свого, аж поки не виросте Шела, син мій. Бо він був подумав: Аби не вмер також він, як брати його. І пішла Тамара, та й осілася в домі батька свого.
GEN|38|12|І минуло багато днів, і вмерла Шуїна дочка, Юдина жінка. А коли Юда був утішений, то пішов до Тімни, до стрижіїв отари своєї, він і Хіра, товариш його адулламітянин.
GEN|38|13|А Тамарі розповіли, кажучи: Ось тесть твій іде до Тімни стригти отару свою.
GEN|38|14|І зняла вона з себе одежу вдівства свого, і покрилася покривалом, і закрилася. І сіла вона при брамі Енаїм, що по дорозі до Тімни. Бо знала вона, що виріс Шела, а вона не віддана йому за жінку.
GEN|38|15|І побачив її Юда, і прийняв її за блудницю, бо закрила вона обличчя своє.
GEN|38|16|І він збочив до неї на дорогу й сказав: А ну но я ввійду до тебе! Бо він не знав, що вона невістка його. А вона відказала: Що даси мені, коли прийдеш до мене?
GEN|38|17|А він відказав: Я пошлю козлятко з отари. І сказала вона: Якщо даси заставу, аж поки пришлеш.
GEN|38|18|А він відказав: Яка та застава, що дам я тобі? Та сказала: Печатка твоя, і шнурок твій, і палиця твоя, що в руці твоїй. І він дав їй, і зійшовся з нею, а вона завагітніла від нього.
GEN|38|19|І встала вона та й пішла, і зняла покривало своє з себе, і зодягнула одежу вдівства свого.
GEN|38|20|А Юда послав козлятко через приятеля свого адулламітянина, щоб узяти заставу з руки тієї жінки. Та він не знайшов її.
GEN|38|21|І запитав він людей її місця, говорячи: Де та блудниця, що була в Енаїм при дорозі? Вони відказали: Не була тут блудниця.
GEN|38|22|І вернувся він до Юди й сказав: Не знайшов я її, а також люди місця того говорили: Не була тут блудниця.
GEN|38|23|І сказав Юда: Нехай візьме собі ту заставу, щоб ми не стали на ганьбу. Ось я послав був те козлятко, та її не знайшов ти.
GEN|38|24|І сталося так десь по трьох місяцях, і розповіджено Юді, говорячи: Упала в блуд Тамара, твоя невістка, і ось завагітніла вона через блуд. А Юда сказав: Виведіть її, і нехай буде спалена.
GEN|38|25|Коли її вивели, то послала вона до тестя свого, говорячи: Я завагітніла від чоловіка, що це належить йому. І сказала: Пізнай но, чия то печатка, і шнури, і ця палиця?
GEN|38|26|І пізнав Юда й сказав: Вона стала справедливіша від мене, бо я не дав її Шелі, синові своєму. І вже більше не знав він її.
GEN|38|27|І сталося в часі, як родила вона, а ось близнята в утробі її.
GEN|38|28|І сталося, як родила вона, показалася рука одного; і взяла баба-сповитуха, і пов'язала на руку йому нитку червону, говорячи: Цей вийшов найперше.
GEN|38|29|І сталося, що він втягнув свою руку, а ось вийшов його брат. І сказала вона: Нащо ти роздер для себе перепону? І назвала ім'я йому Перец.
GEN|38|30|А потім вийшов брат його, що на руці його була нитка червона. І вона назвала ім'я йому: Зерах.
GEN|39|1|А Йосип був відведений до Єгипту. І купив його Потіфар, царедворець фараонів, начальник царської сторожі, муж єгиптянин, з руки ізмаїльтян, що звели його туди.
GEN|39|2|І був Господь з Йосипом, а він став чоловіком, що мав щастя. І пробував він у домі свого пана єгиптянина.
GEN|39|3|І побачив його пан, що Господь з ним, і що в усьому, що він робить, Господь щастить у руці його.
GEN|39|4|І Йосип знайшов милість в очах його, і служив йому. А той призначив його над домом своїм, і все, що мав, віддав в його руку.
GEN|39|5|І сталося, відколи він призначив його в домі своїм, і над усім, що він мав, то поблагословив Господь дім єгиптянина через Йосипа. І було благословення Господнє в усьому, що він мав, у домі й на полі.
GEN|39|6|І він позоставив усе, що мав, у руці Йосиповій. І не знав він при ньому нічого, окрім хліба, що їв. А Йосип був гарного стану та вродливого вигляду.
GEN|39|7|І сталося по тих пригодах, і звела свої очі на Йосипа жінка пана його. І сказала вона: Ляж зо мною!
GEN|39|8|А він відмовився, і сказав до жінки пана свого: Тож пан мій не знає при мені нічого у домі, а все, що його, він дав у мою руку.
GEN|39|9|Нема більшого в цім домі від мене, і він не стримав від мене нічого, хібащо тебе, бо ти жінка його. Як же я вчиню це велике зло, і згрішу перед Богом?
GEN|39|10|І сталося, що вона день-у-день говорила Йосипові, а він не слухав її, щоб лягти при ній і бути з нею.
GEN|39|11|І сталося одного дня, і прийшов він додому робити діло своє, а там у домі не було нікого з людей дому.
GEN|39|12|І схопила вона його за одежу його, кажучи: Лягай же зо мною! А він позоставив свою одежу в її руці, та й утік, і вибіг надвір.
GEN|39|13|І сталося, як побачила вона, що він позоставив свою одежу в її руці та й утік надвір,
GEN|39|14|то покликала людей свого дому, та й сказала їм, говорячи: Дивіться, він припровадив нам якогось єврея, щоб той забавлявся нами! Він прийшов був до мене, щоб покластись зо мною, та я закричала сильним голосом.
GEN|39|15|І сталося, як почув він, що я підняла свій голос і закричала, то позоставив одежу свою в мене, та й утік, і вибіг надвір...
GEN|39|16|І я поклала його одежу при собі аж до приходу пана його до свого дому.
GEN|39|17|І вона переказала йому цими словами, говорячи: До мене прийшов був оцей раб єврей, що ти його привів до нас, щоб забавлятися мною.
GEN|39|18|І сталося, як підняла я свій голос і закричала, то він позоставив свою одежу при мені, та й утік надвір.
GEN|39|19|І сталося, як почув пан його слова своєї жінки, що оповідала йому, кажучи: Отакі то речі вчинив мені твій раб, то запалився гнів його.
GEN|39|20|І взяв його Йосипів пан, та й віддав його до дому в'язничного, до місця, де були ув'язнені царські в'язні. І пробував він там у тім домі в'язничнім.
GEN|39|21|А Господь був із Йосипом, і прихилив до нього милосердя, та дав йому милість в очах начальника в'язничного дому.
GEN|39|22|І начальник в'язничного дому дав у руку Йосипа всіх в'язнів, що були в домі в'язничнім, і все, що там робили, робив він.
GEN|39|23|Начальник в'язничного дому не бачив нічого в руці його, бо Бог був із ним, і що він робив, щастив йому Господь.
GEN|40|1|І сталося по тих пригодах, чашник єгипетського царя та пекар провинилися були панові своєму, цареві єгипетському.
GEN|40|2|І розгнівався фараон на двох своїх евнухів, на начальника чашників і на начальника пекарів.
GEN|40|3|І віддав їх під варту до дому начальника царської сторожі до в'язничного дому, до місця, де Йосип був ув'язнений.
GEN|40|4|А начальник царської сторожі приставив Йосипа до них, і він їм услуговував. І були вони деякий час під вартою.
GEN|40|5|І снився їм обом сон, кожному свій сон, однієї ночі, кожному за значенням його сна, чашникові й пекареві царя єгипетського, що були ув'язнені у в'язничному домі.
GEN|40|6|І прибув до них Йосип уранці, і побачив їх, а вони ось сумні.
GEN|40|7|І запитав він фараонових евнухів, що були з ним під вартою в домі пана його, говорячи: Чого ваші обличчя сьогодні сумні?
GEN|40|8|А вони сказали йому: Снився нам сон, а відгадати його немає кому. І сказав до них Йосип: Чи ж не в Бога відгадки? Розповіджте но мені.
GEN|40|9|І оповів начальник чашників Йосипові свій сон, і сказав йому: Бачив я в сні своїм, ось виноградний кущ передо мною.
GEN|40|10|А в виноградному кущі три виноградні галузки, а він сам ніби розцвів, пустив цвіт, і дозріли грона його ягід.
GEN|40|11|А в моїй руці фараонова чаша. І взяв я ті ягоди, і вичавив їх до фараонової чаші, і дав ту чашу в руку фараона.
GEN|40|12|І сказав йому Йосип: Оце відгадка його: три виноградні галузки це три дні.
GEN|40|13|Ще за три дні підійме фараон твою голову, і верне тебе на твоє становище, і ти даси чашу фараона до руки його за першим звичаєм, як був ти чашником його.
GEN|40|14|Коли ти згадаєш собі про мене, як буде тобі добре, то вчиниш милість мені, коли згадаєш про мене перед фараоном, і випровадиш мене з цього дому.
GEN|40|15|Бо я був справді вкрадений із Краю єврейського, а також тут я не вчинив нічого, щоб мене вкинути до цієї ями.
GEN|40|16|І побачив начальник пекарів, що він добре відгадав, і промовив до Йосипа: І я в сні своїм бачив, ось три коші печива на голові моїй.
GEN|40|17|А в коші горішньому зо всякого пекарського виробу фараонове їдження, а птах їв його з коша з-над моєї голови.
GEN|40|18|І відповів Йосип і сказав: Оце відгадка його: три коші то три дні.
GEN|40|19|Ще за три дні підійме фараон голову твою з тебе, і повісить тебе на дереві, і птах поїсть тіло твоє з тебе.
GEN|40|20|І сталося третього дня, у день народження фараона, і вчинив він гостину для всіх своїх рабів. І підняв він голову начальника чашників і голову начальника пекарів серед своїх рабів.
GEN|40|21|І вернув він начальника чашників на його місце, і він подав чашу в руку фараонову.
GEN|40|22|А начальника пекарів повісив, як відгадав був їм Йосип.
GEN|40|23|Та начальник чашників не пам'ятав про Йосипа, та й забув за нього.
GEN|41|1|І сталося по закінченні двох літ часу, і сниться фараонові, ось він стоїть над Річкою.
GEN|41|2|І ось виходять із Річки семеро корів гарного вигляду й ситого тіла, і паслися на лузі.
GEN|41|3|А ось виходять із Річки за ними семеро корів інших, бридкі виглядом і худі тілом. І вони стали при тих коровах на березі Річки.
GEN|41|4|І корови бридкі виглядом і худі тілом поз'їдали сім корів гарних виглядом і ситих. І прокинувся фараон.
GEN|41|5|І знову заснув він. І снилося йому вдруге, аж ось сходять на однім стеблі семеро колосків здорових та добрих.
GEN|41|6|А ось виростає за ними семеро колосків тонких та спалених східнім вітром.
GEN|41|7|І проковтнули ті тонкі колоски сім колосків здорових та повних. І прокинувся фараон, а то був сон.
GEN|41|8|І сталося рано, і занепокоївся дух його. І послав він, і поскликав усіх ворожбитів Єгипту та всіх мудреців його. І фараон розповів їм свій сон, та ніхто не міг відгадати їх фараонові.
GEN|41|9|І говорив начальник чашників з фараоном, кажучи: Я сьогодні згадую гріхи свої.
GEN|41|10|Розгнівався був фараон на рабів своїх, і вмістив мене під варту дому начальника царської сторожі, мене й начальника пекарів.
GEN|41|11|І однієї ночі снився нам сон, мені та йому, кожному снився сон за своїм значенням.
GEN|41|12|А там з нами був єврейський юнак, раб начальника царської сторожі. І ми розповіли йому, а він відгадав нам наші сни, кожному за сном його відгадав.
GEN|41|13|І сталося, як він відгадав нам, так і трапилося: мене ти вернув на становище моє, а того повісив.
GEN|41|14|І послав фараон, і покликав Йосипа, і його сквапно вивели з в'язниці. І оголився, і змінив одежу свою, і він прибув до фараона.
GEN|41|15|І промовив фараон до Йосипа: Снився мені сон, та нема, хто б відгадав його. А я чув про тебе таке: ти вислухуєш сон, щоб відгадати його.
GEN|41|16|А Йосип сказав до фараона, говорячи: Не я, Бог дасть у відповідь мир фараонові.
GEN|41|17|І сказав фараон до Йосипа: Бачив я в сні своїм ось я стою на березі Річки.
GEN|41|18|І ось виходять із Річки семеро корів ситих тілом і гарних виглядом. І вони паслися на лузі.
GEN|41|19|А ось виходять за ними семеро корів інші, бідні та дуже бридкі виглядом і худі тілом. Таких бридких, як вони, я не бачив у всьому краї єгипетському.
GEN|41|20|І корови худі та бридкі поз'їдали сім корів перших ситих.
GEN|41|21|І ввійшли вони до черева їхнього, та не було знати, що ввійшли вони до черева їхнього, і вигляд їх був лихий, як на початку. І я прокинувся.
GEN|41|22|І побачив я в сні своїм знов, аж ось сходять на однім стеблі семеро колосків повних та добрих.
GEN|41|23|А ось виростає за ними семеро колосків худих, тонких, спалених східнім вітром.
GEN|41|24|І проковтнули ті тонкі колоски сім колосків добрих. І розповів я те ворожбитам, та не було, хто б мені роз'яснив.
GEN|41|25|І сказав Йосип до фараона: Сон фараонів один він. Що Бог робить, те Він звістив фараонові.
GEN|41|26|Семеро корів добрих то сім літ, і семеро колосків добрих сім літ вони. А сон один він.
GEN|41|27|А сім корів худих і бридких, що вийшли за ними, сім літ вони, і сім колосків порожніх і спалених східнім вітром то будуть сім літ голодних.
GEN|41|28|Оце та річ, що я сказав був фараонові: Що Бог робить, те Він показав фараонові.
GEN|41|29|Ось приходять сім літ, великий достаток у всім краї єгипетськім.
GEN|41|30|А по них настануть сім літ голодних, і буде забутий увесь той достаток в єгипетській землі, і голод винищить край.
GEN|41|31|І не буде видно того достатку в краї через той голод, що настане потім, бо він буде дуже тяжкий.
GEN|41|32|А що сон повторився фараонові двічі, це значить, що справа ця постановлена від Бога, і Бог незабаром виконає її.
GEN|41|33|А тепер нехай фараон наздрить чоловіка розумного й мудрого, і нехай поставить його над єгипетською землею.
GEN|41|34|Нехай учинить фараон, і нехай призначить урядників над краєм, і нехай за сім літ достатку збирає п'ятину врожаю єгипетської землі.
GEN|41|35|І нехай вони позбирають усю їжу тих добрих років, що приходять, і нехай вони позбирають збіжжя під руку фараонову, на їжу по містах, і нехай бережуть.
GEN|41|36|І буде та їжа на запас для краю на сім літ голодних, що настануть в єгипетській землі, і край не буде знищений голодом.
GEN|41|37|І була ця річ добра в очах фараона та в очах усіх його рабів.
GEN|41|38|І сказав фараон своїм рабам: Чи знайдеться чоловік, як оцей, що Дух Божий у нім?
GEN|41|39|І сказав фараон Йосипові: Що Бог відкрив тобі це все, то немає такого розумного й мудрого, як ти.
GEN|41|40|Ти будеш над домом моїм, а слів твоїх уст буде слухатися ввесь народ мій. Тільки троном я буду вищий від тебе.
GEN|41|41|І сказав фараон Йосипові: Дивись, я поставив тебе над усім краєм єгипетським.
GEN|41|42|І зняв фараон персня свого з своєї руки, та й дав його на руку Йосипову, і зодягнув його в одежу віссонну, а на шию йому повісив золотого ланцюга.
GEN|41|43|І зробив, що він їздив його другим повозом, і кричали перед обличчям його: Кланяйтеся! І поставив його над усім єгипетським краєм.
GEN|41|44|І сказав фараон Йосипові: Я фараон, а без тебе ніхто не підійме своєї руки та своєї ноги в усім краї єгипетськім.
GEN|41|45|І назвав фараон ім'я Йосипові: Цофнат-Панеах, і дав йому за жінку Оснату, дочку Поті-Фера, жерця Ону. І Йосип піднявся над єгипетським краєм.
GEN|41|46|А Йосип був віку тридцяти літ, коли він став перед лицем фараона, царя єгипетського. І пішов Йосип від лиця фараонового, і перейшов через увесь єгипетський край.
GEN|41|47|А земля в сім літ достатку родила на повні жмені.
GEN|41|48|І зібрав він усю їжу семи літ, що була в єгипетськім краї, і вмістив їжу по містах: їжу поля міста, що навколо нього, вмістив у ньому.
GEN|41|49|І зібрав Йосип збіжжя дуже багато, як морський пісок, аж перестав рахувати, бо не було вже числа.
GEN|41|50|А Йосипові, поки прийшов рік голодний, уродилися два сини, що вродила йому Осната, дочка Поті-Фера, жерця Ону.
GEN|41|51|І назвав Йосип ім'я перворідному: Манасія, бо Бог зробив мені, що я забув усе своє терпіння та ввесь дім мого батька.
GEN|41|52|А ймення другому назвав: Єфрем, бо розмножив мене Бог у краї недолі моєї.
GEN|41|53|І скінчилися сім літ достатку, що були в єгипетськім краї.
GEN|41|54|І зачали наступати сім літ голодні, як сказав був Йосип. І був голод по всіх краях, а в усім єгипетськім краї був хліб.
GEN|41|55|Але виголоднів увесь єгипетський край, а народ став кричати до фараона про хліб. І сказав фараон усьому Єгиптові: Ідіть до Йосипа. Що він вам скаже, те робіть.
GEN|41|56|І був той голод на всій поверхні землі. І відчинив Йосип усе, що було в них, і продавав поживу Єгиптові. А голод зміцнявся в єгипетськім краї.
GEN|41|57|І прибували зо всієї землі до Йосипа купити поживи, бо голод зміцнявся по всій землі.
GEN|42|1|А Яків побачив, що в Єгипті є хліб. І сказав Яків до синів своїх: Пощо ви споглядаєте один на одного?
GEN|42|2|І сказав він: Ось чув я, що в Єгипті є хліб; зійдіть туди, і купіть нам хліба ізвідти, і будемо жити, і не помремо.
GEN|42|3|І зійшли десятеро Йосипових братів купити збіжжя з Єгипту.
GEN|42|4|А Веніямина, Йосипового брата, Яків не послав із братами його, бо сказав: Щоб не спіткало його яке нещастя!
GEN|42|5|І прибули Ізраїлеві сини купити хліба разом з іншими, що приходили, бо був голод у Краї ханаанськім.
GEN|42|6|А Йосип він володар над тим краєм, він продавав хліб усьому народові тієї землі. І прибули Йосипові брати, та й уклонилися йому обличчям до землі.
GEN|42|7|І побачив Йосип братів своїх, і пізнав їх, та не дав пізнати себе. І говорив із ними суворо, і промовив до них: Звідкіля прибули ви? А вони відказали: З ханаанського Краю купити їжі.
GEN|42|8|І пізнав Йосип братів своїх, а вони не впізнали його.
GEN|42|9|І згадав Йосип сни, що про них йому снились були. І сказав він до них: Ви шпигуни! Ви прибули підглянути слабі місця цієї землі.
GEN|42|10|А вони відказали йому: Ні, пане мій, а раби твої прибули купити їжі.
GEN|42|11|Ми всі сини одного чоловіка, ми правдиві. Раби твої не були шпигунами!
GEN|42|12|Він же промовив до них: Ні, бо ви прийшли підглянути слабі місця цієї землі!
GEN|42|13|А вони відказали: Дванадцятеро твоїх рабів брати ми, сини одного чоловіка в ханаанському Краї. А наймолодший тепер із батьком нашим, а одного нема.
GEN|42|14|І промовив їм Йосип: Оце те, що я сказав був до вас, говорячи: Ви шпигуни.
GEN|42|15|Оцим ви будете випробувані: Клянуся життям фараоновим, що ви не вийдете звідси, якщо не прийде сюди наймолодший ваш брат!
GEN|42|16|Пошліть з-поміж себе одного, і нехай візьме вашого брата, а ви будете ув'язнені. І слова ваші будуть піддані пробі, чи правда з вами; а коли ні, клянуся життям фараоновим, що ви шпигуни!
GEN|42|17|І він забрав їх під варту на три дні.
GEN|42|18|А третього дня Йосип промовив до них: Зробіть це і живіть. Я Бога боюся,
GEN|42|19|якщо ви правдиві. Один брат ваш буде ув'язнений в домі вашої варти, а ви йдіть, принесіть хліба для заспокоєння голоду ваших домів.
GEN|42|20|А свого наймолодшого брата приведіть до мене, і будуть потверджені ваші слова, а ви не повмираєте. І вони зробили так.
GEN|42|21|І говорили вони один одному: Справді, винні ми за нашого брата, бо ми бачили недолю душі його, коли він благав нас, а ми не послухали... Тому то прийшло це нещастя на нас!
GEN|42|22|І відповів їм Рувим, говорячи: Чи не говорив я вам, кажучи: Не грішіть проти хлопця, та ви не послухали. А оце й кров його жадається...
GEN|42|23|А вони не знали, що Йосип їх розуміє, бо був поміж ними перекладач.
GEN|42|24|А він відвернувся від них та й заплакав... І вернувся до них, і говорив із ними. І взяв від них Симеона, та й зв'язав його на їхніх очах.
GEN|42|25|А Йосип наказав, щоб наповнили їхні мішки збіжжям, а срібло їхнє вернули кожному до його мішка, і дали їм поживи на дорогу. І їм зроблено так.
GEN|42|26|І понесли вони хліб свій на ослах своїх, і пішли звідти.
GEN|42|27|І відкрив один мішка свого, щоб ослові своєму дати паші на нічлігу, та й побачив срібло своє, а воно ось в отворі мішка його!
GEN|42|28|І сказав він братам своїм: Повернене срібло моє, і ось воно в мішку моїм! І завмерло їм серце, і вони затремтіли, говорячи один до одного: Що це Бог нам зробив?
GEN|42|29|І прибули вони до Якова, батька свого, до Краю ханаанського, і розповіли йому все, що їх спіткало було, говорячи:
GEN|42|30|Той муж, пан того краю, говорив із нами суворо, і прийняв був нас як шпигунів того краю.
GEN|42|31|А ми сказали йому: Ми правдиві, не були ми шпигунами!
GEN|42|32|Ми дванадцятеро братів, сини нашого батька. Одного нема, а наймолодший тепер з нашим батьком у ханаанському Краї.
GEN|42|33|І сказав до нас муж той, пан того краю: З того пізнаю, що правдиві ви, зоставте зо мною одного вашого брата, а на голод домів ваших візьміть хліб та й ідіть.
GEN|42|34|І приведіть до мене брата вашого найменшого, і буду я знати, що ви не шпигуни, що ви правдиві. Тоді віддам вам вашого брата, і ви можете переходити цей край для купівлі.
GEN|42|35|І сталося, вони випорожнювали мішки свої, а ось у кожного вузлик срібла його в його мішку! І побачили вузлики срібла свого, вони та їх батько, і полякались...
GEN|42|36|І сказав до них Яків, їх батько: Ви позбавили мене дітей, Йосипа нема, і Симеона нема, а тепер Веніямина заберете? Усе те на мене!
GEN|42|37|І промовив Рувим до батька свого, кажучи: Двох синів моїх уб'єш, коли не приведу його до тебе! Дай же його на руку мою, а я поверну його до тебе.
GEN|42|38|А той відказав: Не зійде з вами мій син, бо брат його вмер, а він сам позостався... А трапиться йому нещастя в дорозі, якою підете, то в смутку зведете мою сивину до шеолу!...
GEN|43|1|А голод став тяжкий у тім Краї.
GEN|43|2|І сталося, як вони скінчили їсти хліб, що привезли були з Єгипту, то сказав до них батько їх: Верніться, купіть нам трохи їжі!
GEN|43|3|І сказав йому Юда, говорячи: Рішуче освідчив нам той муж, кажучи: Не побачите лиця мого без вашого брата з вами!
GEN|43|4|Як ти пошлеш брата нашого з нами, то ми зійдемо, і купимо тобі їжі.
GEN|43|5|А коли не пошлеш, не зійдемо, бо муж той сказав нам: Не побачите лиця мого без вашого брата з вами.
GEN|43|6|І промовив Ізраїль: Нащо зло ви вчинили мені, що сказали тому мужеві, що ще маєте брата?
GEN|43|7|А вони відказали: Розпитуючи, випитував той муж про нас та про місце нашого народження, говорячи: Чи батько ваш іще живий? Чи є в вас брат? І ми розповіли йому відповідно до цих слів. Чи могли ми знати, що скаже: Приведіть вашого брата?
GEN|43|8|І сказав Юда до Ізраїля, батька свого: Пошли ж цього юнака зо мною, і встаньмо, та й ходім, і будемо жити, і не повмираємо і ми, і ти, і наші діти.
GEN|43|9|Я поручуся за нього, з моєї руки будеш його ти жадати! Коли я не приведу його до тебе, і не поставлю перед лицем твоїм, то буду винним перед тобою по всі дні!
GEN|43|10|А коли б ми були не відтягалися, то тепер уже б вернулися були два рази.
GEN|43|11|І сказав їм Ізраїль, їх батько: Коли так, то зробіть ви оце. Візьміть із плодів цього Краю, і віднесіть дарунка мужеві тому: трохи бальзаму, і трохи меду, пахощів, і ладану, дактилів, і мигдалів.
GEN|43|12|А срібла візьміть удвоє в руку свою. А срібло, повернене в отвір ваших мішків, верніть своєю рукою, може то помилка.
GEN|43|13|А брата вашого заберіть, і встаньте, ідіть до того мужа.
GEN|43|14|А Бог Всемогутній нехай дасть вам милосердя перед лицем того мужа, і нехай він відпустить вам другого вашого брата й Веніямина. А я, певно стратив сина свого!...
GEN|43|15|І взяли ті люди того дарунка, і взяли вдвоє срібла в руку свою, і Веніямина, і встали, та й зійшли до Єгипту. І стали вони перед лицем Йосиповим.
GEN|43|16|І побачив Йосип Веніямина з ними, і сказав до того, що був над його домом: Упровадь цих людей до дому, і нехай заріжуть худобину, і приготуй, бо зо мною будуть їсти ці люди опівдні.
GEN|43|17|І той чоловік зробив, як Йосип сказав був. І впровадив той чоловік тих людей до Йосипового дому.
GEN|43|18|І полякалися ті люди, що були впроваджені до Йосипового дому. І сказали вони: Через срібло, повернене напочатку в наших мішках, ми впроваджені, щоб причепитись до нас, і напасти на нас, і забрати за рабів нас та наші осли...
GEN|43|19|І приступили вони до чоловіка, що над домом Йосиповим, та й говорили до нього при вході в дім.
GEN|43|20|І сказали вони: Послухай, о пане мій, ми зійшли були напочатку купити їжі.
GEN|43|21|І сталося, коли ми прийшли на нічліг, і відкрили мішки свої, а ось срібло кожного в отворі мішка його, наше срібло за вагою його! І ми вертаємо його нашою рукою!
GEN|43|22|А на купівлю їжі ми знесли нашою рукою інше срібло. Ми не знаємо, хто поклав був наше срібло до наших мішків...
GEN|43|23|А той відказав: Мир вам! Не бійтеся! Бог ваш і Бог вашого батька дав вам скарб до ваших мішків. Срібло ваше прийшло до мене. І вивів до них Симеона.
GEN|43|24|І впровадив той чоловік тих людей до Йосипового дому, і дав води, а вони вмили ноги свої, і дав паші їхнім ослам.
GEN|43|25|І вони приготовили дарунки до приходу Йосипа опівдні, бо почули, що там вони їстимуть хліб.
GEN|43|26|І ввійшов Йосип до дому, а вони принесли йому до дому дарунка, що в їхній руці. І вони поклонилися йому до землі.
GEN|43|27|А він запитав їх про мир і сказав: Чи гаразд вашому батькові старому, про якого ви розповідали? Чи він ще живий?
GEN|43|28|А вони відказали: Гаразд рабові твоєму, батькові нашому. Ще він живий. І вони схилилися, і вклонилися до землі.
GEN|43|29|І звів він очі свої, та й побачив Веніямина, свого брата, сина матері своєї, і промовив: Чи то ваш наймолодший брат, що ви мені розповідали? І сказав: Нехай Бог буде милостивий до тебе, мій сину!
GEN|43|30|І Йосип поспішив, бо порушилася його любов до брата його, і хотів він заплакати. І ввійшов він до іншої кімнати, і заплакав там...
GEN|43|31|І вмив він лице своє, і вийшов, і стримався, та й сказав: Покладіть хліба!
GEN|43|32|І поклали йому окремо, а їм окремо, й єгиптянам, що їли з ним, окремо, бо єгиптяни не можуть їсти хліб з євреями, бо це огида для Єгипту.
GEN|43|33|І вони посідали перед ним, перворідний за перворідством своїм, а молодший за молодістю своєю. І здивувалися ці люди один перед одним.
GEN|43|34|І він посилав дари страви від себе до них. А дар Веніяминів був більший від дару всіх їх уп'ятеро. І пили вони, і повпивалися з ним.
GEN|44|1|І наказав він тому, що над домом його, говорячи: Понаповнюй мішки цих людей їжею, скільки зможуть вони нести. І поклади срібло кожного до отвору мішка його.
GEN|44|2|А чашу мою, чашу срібну, поклади до отвору мішка наймолодшого, та срібло за хліб його. І зробив той за словом Йосиповим, яке він сказав був.
GEN|44|3|Розвиднилось рано вранці, і люди ці були відпущені, вони та їхні осли.
GEN|44|4|Вони вийшли з міста, ще не віддалилися, а Йосип сказав до того, що над домом його: Устань, побіжи за тими людьми, і дожени їх, та й скажи їм: Нащо ви заплатили злом за добро?
GEN|44|5|Хіба це не та чаша, що з неї п'є пан мій, і він, ворожачи, ворожить нею? І зле ви зробили, що вчинили таке.
GEN|44|6|І той їх догнав, і сказав їм ті слова.
GEN|44|7|А вони відказали йому: Нащо пан мій говорить отакі то слова? Далеке рабам твоїм, щоб зробити таку річ...
GEN|44|8|Таж срібло, що знайшли ми в отворах наших мішків, ми вернули тобі з Краю ханаанського. А як би ми вкрали з дому пана твого срібло чи золото?
GEN|44|9|У кого із рабів твоїх вона, чаша, буде знайдена, то помре він, а також ми станемо рабами моєму панові.
GEN|44|10|А той відказав: Тож тепер, як ви сказали, так нехай буде воно! У кого вона знайдена буде, той стане мені за раба, а ви будете чисті.
GEN|44|11|І поспішно поспускали вони кожен свого мішка на землю. І порозв'язували кожен мішка свого.
GEN|44|12|І став він шукати. Розпочав від найстаршого, а скінчив наймолодшим. І знайдена чаша в мішку Веніяминовім!
GEN|44|13|І пороздирали вони свою одіж!... І кожен нав'ючив осла свого, і вернулись до міста.
GEN|44|14|І ввійшли Юда й брати його до дому Йосипа, а він ще був там. І попадали вони перед лицем його на землю.
GEN|44|15|І сказав до них Йосип: Що це за вчинок, що ви зробили? Хіба ви не знали, що справді відгадає такий муж, як я?
GEN|44|16|А Юда промовив: Що ми скажемо панові моєму? Що будемо говорити? Чим виправдаємось? Бог знайшов провину твоїх рабів! Ось ми раби панові моєму, і ми, і той, що в руці його була знайдена чаша.
GEN|44|17|А Йосип відказав: Далеке мені, щоб зробити оце. Чоловік, що в руці його була знайдена чаша, він буде мені за раба! А ви йдіть із миром до вашого батька.
GEN|44|18|І приступив до нього Юда та й промовив: О мій пане, нехай скаже раб твій слово до ушей пана свого, і нехай не палає гнів твій на раба твого, бо ти такий, як фараон.
GEN|44|19|Пан мій запитав був рабів своїх, говорячи: Чи є в вас батько або брат?
GEN|44|20|І сказали ми до пана мого: Є в нас батько старий та мале дитя його старости, а брат його вмер. І позостався він сам у своєї матері, а батько його любить.
GEN|44|21|А ти був сказав своїм рабам: Зведіть до мене його, і нехай я кину своїм оком на нього.
GEN|44|22|І сказали ми до пана мого: Не може той хлопець покинути батька свого. А покине він батька свого, то помре той.
GEN|44|23|А ти сказав своїм рабам: Коли не зійде з вами наймолодший ваш брат, не побачите більше лиця мого.
GEN|44|24|І сталося, коли ми зійшли були до раба твого, до нашого батька, то ми розповіли йому слова мого пана.
GEN|44|25|А батько наш сказав: Верніться, купіть нам трохи їжі.
GEN|44|26|А ми відказали: Не можемо зійти.
GEN|44|27|І сказав до нас раб твій, наш батько: Ви знаєте, що двох була породила мені жінка моя.
GEN|44|28|Та пішов від мене один, і я сказав: справді, дійсно розшарпаний він... І я не бачив його аж дотепер.
GEN|44|29|А заберете ви також цього від мене, і спіткає його нещастя, то зведете ви сивину мою цим злом до шеолу.
GEN|44|30|А тепер, коли я прийду до раба твого, мого батька, а юнака не буде з нами, а душа його зв'язана з душею тією,
GEN|44|31|То станеться, коли він побачить, що юнака нема, то помре. І зведуть твої раби сивину раба твого, нашого батька, у смутку до шеолу...
GEN|44|32|Бо раб твій поручився за юнака батькові своєму, кажучи: Коли я не приведу його до тебе, то згрішу перед батьком своїм на всі дні!
GEN|44|33|А тепер нехай же сяде твій раб замість того юнака за раба панові моєму. А юнак нехай іде з своїми братами!...
GEN|44|34|Бо як я прийду до батька свого, а юнака зо мною нема? Щоб не побачити мені того нещастя, що спіткає мого батька.
GEN|45|1|І не міг Йосип здержатися при всіх, що стояли біля нього, та й закричав: Виведіть усіх людей від мене! І не було з ним нікого, коли Йосип відкрився браттям своїм.
GEN|45|2|І він голосно заплакав, і почули єгиптяни, і почув дім фараонів.
GEN|45|3|І Йосип промовив до браттів своїх: Я Йосип... Чи живий ще мій батько?... І не могли його браття йому відповісти, бо вони налякались його...
GEN|45|4|А Йосип промовив до братів своїх: Підійдіть же до мене! І вони підійшли, а він проказав: Я Йосип, ваш брат, якого ви продали були до Єгипту...
GEN|45|5|А тепер не сумуйте, і нехай не буде жалю в ваших очах, що ви продали мене сюди, бо то Бог послав мене перед вами для виживлення.
GEN|45|6|Бо ось два роки голод на землі, і ще буде п'ять літ, що не буде орки та жнив.
GEN|45|7|І послав мене Бог перед вами зробити для вас, щоб ви позостались на землі, і щоб утримати для вас при житті велике число спасених.
GEN|45|8|І виходить тепер, не ви послали мене сюди, але Бог. І Він зробив мене батьком фараоновим і паном усього дому його, і володарем усього краю єгипетського.
GEN|45|9|Поспішіть, і йдіть до батька мого, та й скажіть йому: Отак сказав син твій Йосип: Бог зробив мене володарем усього Єгипту. Зійди ж до мене, не гайся.
GEN|45|10|І осядь у землі Ґошен, і будеш близький до мене ти, і сини твої, і сини синів твоїх, і дрібна та велика худоба твоя, і все, що твоє.
GEN|45|11|І прогодую тебе там, бо голод буде ще п'ять років, щоб не збіднів ти, і дім твій, і все, що твоє.
GEN|45|12|І ось очі ваші й очі брата мого Веніямина бачать, що це мої уста говорять до вас.
GEN|45|13|І оповісте батькові моєму про всю славу мою в Єгипті, та про все, що ви бачили. І поспішіть, і приведіть вашого батька сюди.
GEN|45|14|І впав він на шию Веніямину, братові своєму, та й заплакав, і Веніямин плакав на шиї його...
GEN|45|15|І цілував він усіх братів своїх, і плакав над ними... А потому говорили брати його з ним.
GEN|45|16|І розголошено в домі фараоновім чутку, говорячи: Прийшли Йосипові брати! І було це добре в очах фараонових та в очах його рабів.
GEN|45|17|І промовив фараон до Йосипа: Скажи своїм братам: Зробіть оце: Понав'ючуйте худобу свою, та й ідіть, прибудьте до Краю ханаанського.
GEN|45|18|І заберіть вашого батька й доми ваші, та й прийдіть до мене, а я дам вам добра єгипетського краю. І споживайте ситість землі.
GEN|45|19|А ти одержав наказа сказати: Зробіть це: Візьміть собі з єгипетського краю вози для ваших дітей та для ваших жінок, і привезіть свого батька й прибудьте.
GEN|45|20|А око ваше нехай не жалує ваших речей, бо добро всього єгипетського краю ваше воно.
GEN|45|21|І зробили так Ізраїлеві сини. А Йосип дав їм вози на приказ фараонів, і дав їм поживи на дорогу.
GEN|45|22|І дав усім їм кожному переміни одежі, а Веніяминові дав три сотні срібла та п'ять перемін одежі.
GEN|45|23|А батькові своєму послав він оце: десять ослів, нав'ючених з добра Єгипту, і десять ослиць, нав'ючених збіжжям, і хліб, і поживу для батька його на дорогу.
GEN|45|24|І відпустив він своїх братів, і вони пішли. І сказав він до них: Не сваріться в дорозі!
GEN|45|25|І вийшли вони з Єгипту, та й прибули до ханаанського Краю, до Якова, батька свого.
GEN|45|26|І розповіли йому, кажучи: Ще Йосип живий, і що він панує над усім єгипетським краєм. І зомліло серце його, бо він не повірив був їм...
GEN|45|27|І переказували йому всі слова Йосипові, що говорив він до них. І як побачив він вози, що послав Йосип, щоб везти його, то ожив дух Якова, їхнього батька.
GEN|45|28|І промовив Ізраїль: Досить! Ще живий Йосип, мій син! Піду ж та побачу його, поки помру!
GEN|46|1|І вирушив Ізраїль, і все, що його, і прибув до Беер-Шеви, і приніс жертви Богові батька свого Ісака.
GEN|46|2|І промовив Бог до Ізраїля в нічному видінні, і сказав: Якове, Якове! А той відказав: Ось я!
GEN|46|3|І сказав Він: Я Той Бог, Бог батька твого. Не бійся зійти до Єгипту, бо Я вчиню тебе там великим народом.
GEN|46|4|Я зійду з тобою до Єгипту, і Я також, виводячи, виведу тебе, а Йосип закриє рукою своєю очі твої.
GEN|46|5|І встав Яків з Беер-Шеви. І повезли Ізраїлеві сини свого батька Якова, і дітей своїх, і жінок своїх возами, що послав фараон, щоб привезти його.
GEN|46|6|І взяли вони стада свої, і маєток свій, що набули в землі ханаанській, і прибули до Єгипту Яків та ввесь рід його з ним.
GEN|46|7|Він привів із собою до Єгипту синів своїх, і синів своїх синів з собою, дочок своїх, і дочок синів своїх, і ввесь рід свій.
GEN|46|8|А оце ймення синів Ізраїлевих, що прибули до Єгипту: Яків та сини його: перворідний Яковів Рувим.
GEN|46|9|І сини Рувимові: Ханох, і Паллу, і Хецрон, і Кармі.
GEN|46|10|І сини Симеонові: Ємуїл, і Ямін, і Огад, і Яхін, і Цохар, і Саул, син ханаанеянки.
GEN|46|11|І сини Левієві: Ґершон, Кегат і Мерарі.
GEN|46|12|І сини Юдині: Ер, і Онан, і Шела, і Перец, і Зерах. І вмер Ер і Онан у ханаанській землі. А сини Перецеві були: Хецрон і Хамул.
GEN|46|13|І сини Іссахарові: Тола, і Цувва, і Йов, і Шимрон.
GEN|46|14|І сини Завулонові: Серед, і Елон, і Яхлеїл.
GEN|46|15|Оце сини Ліїні, що вродила вона Якову в Падані арамейськім, та дочку його Діну. Усіх душ синів його й дочок його тридцять три.
GEN|46|16|І сини Ґадові: Ціфйон, і Хаґґі, Шуні, і Ецбон, Ері, і Ароді, і Ар'їлі.
GEN|46|17|І сини Асирові: Їмна, і Їшва, і Їшві, і Верія, і Сірах, сестра їх. І сини Верії: Хевер і Малкіїл.
GEN|46|18|Оце сини Зілпи, що Лаван був дав її своїй дочці Лії, а вона вродила їх Якову, шістнадцять душ.
GEN|46|19|Сини Рахілі, жінки Якова: Йосип і Веніямин.
GEN|46|20|І вродилися Йосипові в єгипетськім краї Манасія та Єфрем, що їх уродила йому Оснат, дочка Поті-Фера, жерця Ону.
GEN|46|21|І сини Веніяминові: Бела, і Бехер, і Ашбел, Ґера, і Нааман, Ехі, і Рош, Муппім, і Хуппім, і Ард.
GEN|46|22|Оце сини Рахілині, що вродилися Якову, усіх душ чотирнадцять.
GEN|46|23|І сини Данові: Хушім.
GEN|46|24|І сини Нефталимові: Яхсеїл, і Ґуні, і Єцер, і Шіллем.
GEN|46|25|Оце сини Білги, що її Лаван дав був своїй дочці Рахілі. І вона породила їх Якову, усіх душ сім.
GEN|46|26|Усіх душ, що прийшли з Яковом в Єгипет, що походять із стегон його, окрім жінок синів Якова, усіх душ шістдесят і шість.
GEN|46|27|А сини Йосипа, що народилися йому в Єгипті, дві душі. Усіх душ дому Якова, що прийшли були до Єгипту, сімдесят.
GEN|46|28|І послав він перед собою Юду до Йосипа, щоб показував перед ним дорогу до Ґошену. І прибули вони до краю Ґошен.
GEN|46|29|І запріг Йосип свою колесницю, і вирушив назустріч батькові своєму Ізраїлеві до Ґошену. І він показався йому, і впав йому на шию, та й плакав довго на шиї його...
GEN|46|30|І промовив Ізраїль до Йосипа: Нехай тепер помру я, побачивши обличчя твоє, що ти ще живий!
GEN|46|31|А Йосип промовив до своїх братів і до дому батька свого: Піду й розкажу фараонові, та й повім йому: Брати мої й дім батька мого, що були в Краї ханаанськім, прибули до мене.
GEN|46|32|А люди ці пастухи отари, бо були скотарі. І вони припровадили дрібну та велику худобу свою, і все, що їхнє було.
GEN|46|33|І станеться, коли покличе вас фараон і скаже: Яке ваше зайняття?
GEN|46|34|то ви відкажете: Скотарями були твої раби від молодости своєї аж дотепер, і ми, і батьки наші, щоб ви осіли в країні Ґошен, бо для Єгипту кожен пастух отари огида.
GEN|47|1|І прийшов Йосип, і розповів фараонові та й сказав: Мій батько, і брати мої, і їхні отари, і худоба їх, і все їхнє прибули з ханаанського Краю. І ось вони в країні Ґошен.
GEN|47|2|І взяв він із своїх братів п'ятеро чоловіка, та й поставив їх перед лицем фараоновим.
GEN|47|3|І сказав фараон до братів його: Яке ваше зайняття? А вони відказали фараонові: Пастухи отари раби твої, і ми, і наші батьки.
GEN|47|4|І сказали вони фараонові: Ми прибули, щоб мешкати в краї цім, нема бо паші для отари, що є в рабів твоїх, бо в ханаанському Краї тяжкий голод. А тепер нехай же осядуть раби твої в країні Ґошен.
GEN|47|5|І промовив фараон до Йосипа, говорячи: Батько твій та брати твої прибули до тебе.
GEN|47|6|Єгипетьський край він перед лицем твоїм. У найліпшім місці цього краю осади батька свого та братів своїх, нехай осядуть у країні Ґошен. А коли знаєш, і між ними є здатні люди, то зроби їх зверхниками моєї череди.
GEN|47|7|І привів Йосип батька свого Якова, та й поставив його перед лицем фараоновим. І Яків поблагословив фараона.
GEN|47|8|І промовив фараон до Якова: Скільки днів часу життя твого?
GEN|47|9|А Яків сказав до фараона: Днів часу мандрівки моєї сто й тридцять літ. Короткі та лихі були дні часу життя мого, і не досягли вони днів часу життя батьків моїх у днях часу мандрівки їхньої.
GEN|47|10|І Яків поблагословив фараона, та й вийшов від обличчя фараонового.
GEN|47|11|І осадив Йосип батька свого та братів своїх, і дав їм володіння в єгипетській країні, у найкращім місці цієї землі у країні Рамесес, як наказав був фараон.
GEN|47|12|І постачав Йосип хліб для батька свого й братів своїх, та для всього дому свого батька відповідно до числа дітей.
GEN|47|13|А хліба не було в усім тім краї, бо голод став дуже тяжкий. І виснажився єгипетський край та Край ханаанський через той голод.
GEN|47|14|І зібрав Йосип усе срібло, що знаходилося в єгипетськім краї та в Краї ханаанськім, за поживу, що вони купували. І Йосип вніс те срібло до фараонового дому.
GEN|47|15|І вичерпалося срібло в краї єгипетськім та в Краї ханаанськім. І прибув увесь Єгипет до Йосипа, говорячи: Дай же нам хліба! Нащо нам умирати перед тобою, тому що вичерпалося срібло?
GEN|47|16|А Йосип сказав: Дайте свою худобу, а я дам вам за худобу вашу, коли вичерпалося срібло.
GEN|47|17|І вони припровадили худобу свою до Йосипа. І дав їм Йосип хліба за коні, і за отари, і за череди худоби, і за осли. І він того року постачав їм хліб за всю їхню худобу.
GEN|47|18|І скінчився той рік, і вони прибули до нього другого року, та й сказали йому: Не скажемо неправди перед паном своїм, що вичерпалося срібло, а череди здобутку в нашого пана. Нічого не зосталося перед нашим паном, хібащо наше тіло та наша земля!
GEN|47|19|Нащо ми маємо вмирати на очах твоїх, і ми, і наша земля? Купи нас та нашу землю за хліб, і будемо ми та наша земля рабами фараонові. А ти дай насіння, і будемо жити, і не помремо, а земля не опустіє...
GEN|47|20|І Йосип купив усю землю єгипетську для фараона, бо єгиптяни спродували кожен поле своє, посилився бо був голод між ними. І стала земля фараоновою.
GEN|47|21|А народ він перепроваджував його до міст від кінця границі Єгипту й аж до кінця її.
GEN|47|22|Тільки землі жерців не купив він, бо для жерців була устава жити на прибутки від фараона. І вони їли свій пай, що давав їм фараон, тому не продали своєї землі.
GEN|47|23|І сказав Йосип до народу: Оце купив я сьогодні для фараона вас і землю вашу. Ось вам насіння, і засійте землю.
GEN|47|24|А настануть жнива, то дасте п'яту частину фараонові, а чотири частині будуть вам на насіння для поля й на їжу вам та тим, хто в домах ваших, та на їжу для ваших дітей.
GEN|47|25|А вони відказали: Ти нас удержав при житті. Нехай же знайдемо милість в очах свого пана, і станемо рабами фараонові.
GEN|47|26|А Йосип поклав це за постанову на єгипетську землю аж до сьогоднішнього дня: на п'яту частину для фараона. Сама тільки земля жерців не стала фараоновою.
GEN|47|27|І осів Ізраїль в єгипетськім краї в країні Ґошен, і набули в нім володіння. І вони розродилися й сильно розмножилися.
GEN|47|28|І жив Яків в єгипетськім краї сімнадцять літ. І були дні Якова, літа життя його, сто літ і сорок і сім літ.
GEN|47|29|І наблизилися дні Ізраїля до смерти. І кликнув він до сина свого до Йосипа, та й промовив йому: Коли знайшов я милість в очах твоїх, поклади руку свою під стегно моє, і вчини зо мною милість та правду: Не поховай мене в Єгипті!
GEN|47|30|І ляжу я з батьками своїми, і ти винесеш мене з Єгипту, і поховаєш мене в їхньому гробі. А той відказав: Я вчиню за словом твоїм.
GEN|47|31|А Яків сказав: Присягни ж мені! І він присягнув йому. І вклонився Ізраїль на зголов'я постелі.
GEN|48|1|І сталося по тих випадках, і сказано було Йосипові: Ось батько твій хворіє. І він узяв із собою обох своїх синів, Манасію та Єфрема.
GEN|48|2|І промовив він до Якова й сказав: Ось до тебе прийшов твій син Йосип! І зміцнився Ізраїль, та й сів на постелі.
GEN|48|3|І сказав Яків до Йосипа: Бог Всемогутній явився був мені в Лузі в землі ханаанській, і поблагословив мене.
GEN|48|4|І сказав Він до мене: Ось Я розплоджу тебе й розмножу тебе, і вчиню тебе громадою народів. А цю землю Я дам нащадкам твоїм по тобі володінням навіки.
GEN|48|5|А тепер два сини твої, уроджені тобі в єгипетськім краї до прибуття мого до тебе до Єгипту, вони мої! Єфрем і Манасія, як Рувим і Симеон, будуть мої.
GEN|48|6|А нащадки твої, що породиш по них, вони будуть твої. Вони будуть зватися на ймення своїх братів у наслідді своїм.
GEN|48|7|А я, коли я прийшов був з Падану, померла мені Рахіль у Краї ханаанськім на дорозі, коли була ще ківра землі, щоб прийти до Ефрати. І я поховав був її там, на дорозі до Ефрати, це Віфлеєм.
GEN|48|8|А Ізраїль побачив синів Йосипових та й сказав: Хто вони?
GEN|48|9|І сказав Йосип до батька свого: Вони мої сини, що Бог дав мені тут. А той відказав: Візьми ж їх до мене, і я їх поблагословлю.
GEN|48|10|А очі Ізраїлеві стали тяжкі від старости, він не міг дивитися. І Йосип підвів їх до нього, а той поцілував їх і пригорнув їх.
GEN|48|11|І сказав Ізраїль до Йосипа: Не сподівався я побачити обличчя твого, а ось Бог дав мені побачити й насіння твоє.
GEN|48|12|І Йосип відвів їх від колін його, та й упав на обличчя своє до землі.
GEN|48|13|І Йосип узяв їх обох, Єфрема своєю правицею від лівиці Ізраїля, а Манасію своєю лівицею від правиці Ізраїля, та й до нього підвів.
GEN|48|14|І простяг Ізраїль правицю свою та й поклав на голову Єфрема, а він молодший, а лівицю свою на голову Манасії. Він схрестив свої руки, хоч Манасія перворідний.
GEN|48|15|І він поблагословив Йосипа, та й промовив: Бог, що перед обличчям Його ходили батьки мої Авраам та Ісак, що пасе мене, відколи існую аж до цього дня,
GEN|48|16|Ангол, що рятує мене від усього лихого, нехай поблагословить цих юнаків, і нехай буде зване в них ім'я моє й ім'я батьків моїх Авраама та Ісака, і нехай вони множаться, як та риба, посеред землі.
GEN|48|17|А Йосип побачив, що батько його кладе правицю свою на голову Єфремову, і було це не до вподоби йому. І він підпер руку батька свого, щоб зняти її з-над голови Єфрема на голову Манасіїну.
GEN|48|18|І сказав Йосип до батька свого: Не так, батьку мій, бо оцей перворідний, поклади правицю свою на його голову!
GEN|48|19|А батько його не хотів, і сказав: Знаю, мій сину, знаю! І він буде народом, і він буде великий, але його менший брат буде більший від нього, а потомство його стане повнею народів.
GEN|48|20|І він поблагословив їх того дня, кажучи: Тобою буде благословляти Ізраїль, говорячи: Нехай Бог учинить тебе як Єфрема і як Манасію! І поставив Єфрема перед Манасією.
GEN|48|21|І сказав Ізраїль до Йосипа: Ось я вмираю... А Бог буде з вами, і поверне вас до Краю ваших батьків!
GEN|48|22|А я тобі дав понад братів твоїх одну частку, яку я взяв був з руки амореянина своїм мечем та луком своїм.
GEN|49|1|І покликав Яків усіх синів своїх та й промовив: Зберіться, а я сповіщу вам, що вас спіткає наприкінці днів.
GEN|49|2|Зійдіться та слухайте ви, сини Якова, і прислухайтеся до Ізраїля, вашого батька!
GEN|49|3|Рувиме, ти мій перворідний, моя міць і початок ти сили моєї, верх величности й верх ти могутности!
GEN|49|4|Ти пінився був, як вода, та не втримаєшся, бо ти увійшов був на ложе свойого отця, і збезчестив його, на постелю мою ти піднявся!
GEN|49|5|Симеон і Левій то брати, їхня зброя знаряддя насильства.
GEN|49|6|Хай до їхньої змови не входить душа моя, і нехай не прилучиться слава моя до їх зборів, бо вони в своїм гніві людину забили, а в своїй самоволі вола копит позбавили...
GEN|49|7|Проклятий гнів їхній, бо сильний, та їхня лютість, тяжка бо вона! Поділю їх я в Якові, і їх розпорошу в Ізраїлі!
GEN|49|8|О Юдо, похвалять тебе твої браття! Рука твоя на шиї твоїх ворогів, сини батька твого тобі вклоняться.
GEN|49|9|Юда лев молодий! Ти, мій сину, вертаєшся з здобичі: прихиливсь він, поклався як лев й як левиця, зведе хто його?
GEN|49|10|Не відійметься берло від Юди, ані з його стегон законодавець, аж прийде Примиритель, що Йому буде послух народів.
GEN|49|11|Він прив'язує до винограду свого молодого осла, а до вибраної виноградини сина ослиці своєї. Він одежу свою буде прати в вині, а шату свою в виноградній крові!
GEN|49|12|Від вина він зробивсь мутноокий, а від молока білозубий.
GEN|49|13|Завулон буде мешкать над берегом морським, над берегом тим, де стають кораблі, а границя його до Сидону.
GEN|49|14|Іссахар то костистий осел, що лежить між кошарами.
GEN|49|15|І побачив він спокій, що добрий, та землю, що стала приємна, і він нахилив свої плечі, щоб нести, і став працювать на податок.
GEN|49|16|Дан буде судить свій народ, як один із Ізраїльських родів.
GEN|49|17|Дан буде вужем при дорозі, змією отруйливою при шляху, що п'яти коневі кусає, і його верхівець позад себе впаде.
GEN|49|18|Спасіння від Тебе чекаю, о Господи!
GEN|49|19|Ґад на нього юрба нападатиме, та він нападе на їх п'яти.
GEN|49|20|Асир його хліб буде ситий, і він буде давати присмаки царські.
GEN|49|21|Нефталим вільна ланя, він прекрасні слова видає.
GEN|49|22|Йосип вітка родюча, вітка родючая над джерелом, її віття по муру спинається.
GEN|49|23|І огірчили його та з луку стріляли, і зненавиділи були стрільці його.
GEN|49|24|Та зостався міцним його лук, і стали пружні рамена його рук, від рук Сильного Якового, звідти Пастир, Твердиня синів Ізраїлевих.
GEN|49|25|Проси ти від Бога, свойого Отця, і Він допоможе тобі, і проси Всемогутнього і Він благословить тебе благословенням небес, що на висоті, благословенням безодні, що долі лежить, благословеннями перс та утроби.
GEN|49|26|Благословення батька твого стали сильніші від благословення батьків моїх, аж до пожаданих висот віковічних. Нехай вони будуть на голову Йосипову, на маківку вибраного з-поміж братів своїх!
GEN|49|27|Веніямин хижий вовк: вранці їсть він ловитву, а на вечір розділює здобич.
GEN|49|28|Оце всі дванадцять племен Ізраїлевих, і те, що говорив їм батько їх. І він поблагословив їх, кожного за благословенням його поблагословив їх.
GEN|49|29|І він наказав їм, і промовив до них: Я прилучаюся до своєї рідні... Поховайте мене при батьках моїх у печері, що на полі Ефрона хіттеянина,
GEN|49|30|у тій печері, що на полі Махпели, що навпроти Мамре в ханаанській землі, яке поле купив був Авраам від Ефрона хіттеянина на володіння для гробу.
GEN|49|31|Там поховано Авраама й жінку його Сарру, там поховали Ісака та його жінку Ревеку, і там поховав я Лію.
GEN|49|32|Поле й печера, що на нім, то добуток від синів Хета.
GEN|49|33|І закінчив Яків заповіта синам своїм, і втягнув свої ноги до ліжка, та й спочив. І він прилучився до своєї рідні.
GEN|50|1|І впав Йосип на лице батька свого, та й плакав над ним, і цілував його.
GEN|50|2|І звелів Йосип рабам своїм лікарям забальзамувати батька його. І забальзамували ці лікарі Ізраїля.
GEN|50|3|І сповнилося йому сорок день, бо так сповняються дні бальзамування. І оплакував його Єгипет сімдесят день.
GEN|50|4|А як минули дні оплакування його, то сказав Йосип до дому фараонового, говорячи: Коли знайшов я ласку в очах ваших, то говоріть до ушей фараонових так:
GEN|50|5|Батько мій заприсяг був мене, говорячи: Ось я вмираю. У гробі моїм, що я собі викопав у Країні ханаанській, там поховаєш мене. А тепер нехай я піду, і поховаю батька свого, та й вернуся.
GEN|50|6|І сказав фараон: Піди, і поховай свого батька, як заприсяг він тебе.
GEN|50|7|І пішов Йосип поховати батька свого, а з ним пішли всі раби фараонові, старші дому його, і всі старші єгипетського краю,
GEN|50|8|і ввесь дім Йосипів, і браття його, і дім батька його. Тільки дітей своїх та дрібну й велику худобу свою вони позоставили в країні Ґошен.
GEN|50|9|І вирушили з ним також колесниці та комонники. І був табір їх дуже великий.
GEN|50|10|І прийшли вони до Ґорен-Атаду, що по другім боці Йордану, і плакали там великим та дуже ревним плачем... І він учинив батькові своєму семиденну жалобу.
GEN|50|11|І побачили мешканці того Краю, ханаанеяни, жалобу в Ґорен-Атаді, та й сказали:
GEN|50|12|І вчинили йому сини його так, як він їм заповів був.
GEN|50|13|І понесли його сини його до ханаанського Краю, та й поховали його в печері поля Махпели, яке поле купив був Авраам на володіння для гробу від хіттеянина Ефрона, навпроти Мамре.
GEN|50|14|А Йосип, як поховав він батька свого, вернувся до Єгипту, він і брати його, та всі, хто ходив з ним ховати батька його.
GEN|50|15|І побачили Йосипові брати, що вмер їхній батько, та й сказали: А що як зненавидить нас Йосип, і справді верне нам усе зло, що ми йому були заподіяли?
GEN|50|16|І переказали вони Йосипові, говорячи: Батько твій заповів був перед своєю смертю, кажучи:
GEN|50|17|Отак скажіть Йосипові: Прошу, вибач гріх братів твоїх та їхню провину, бо вони тобі зло були заподіяли! А тепер вибач гріх рабам Бога батька твого! І заплакав Йосип, як вони говорили до нього...
GEN|50|18|І пішли також браття його, і впали перед лицем його, та й сказали: Ось ми тобі за рабів!
GEN|50|19|А Йосип промовив до них: Не бійтеся, бо хіба ж я замість Бога?
GEN|50|20|Ви задумували були на мене зло, та Бог задумав те на добре, щоб зробити, як вийшло сьогодні, щоб заховати при житті великий народ!
GEN|50|21|А тепер не лякайтеся, я буду утримувати вас та дітей ваших! І він потішав їх, і промовляв до їхнього серця.
GEN|50|22|І осівся Йосип в Єгипті, він та дім батька його. І жив Йосип сто і десять літ.
GEN|50|23|І побачив Йосип в Єфрема дітей третього покоління. Також сини Махіра, сина Манасіїного, були народилися на Йосипові коліна.
GEN|50|24|І сказав Йосип до братів своїх: Я вмираю, а Бог конче згадає вас, і виведе вас із цієї землі до Краю, якого присягнув був Авраамові, Ісакові та Якову.
GEN|50|25|І Йосип заприсяг Ізраїлевих синів, говорячи: Конче згадає Бог вас, а ви винесете звідси кості мої!
GEN|50|26|І впокоївся Йосип у віці ста й десяти літ. І забальзамували його, і він був покладений у труну в Єгипті.
