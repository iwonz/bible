ZEPH|1|1|The word of the LORD that came to Zephaniah the son of Cushi, son of Gedaliah, son of Amariah, son of Hezekiah, in the days of Josiah the son of Amon, king of Judah.
ZEPH|1|2|"I will utterly sweep away everything from the face of the earth," declares the LORD.
ZEPH|1|3|"I will sweep away man and beast; I will sweep away the birds of the heavens and the fish of the sea, and the rubble with the wicked. I will cut off mankind from the face of the earth," declares the LORD.
ZEPH|1|4|"I will stretch out my hand against Judah and against all the inhabitants of Jerusalem; and I will cut off from this place the remnant of Baal and the name of the idolatrous priests along with the priests,
ZEPH|1|5|those who bow down on the roofs to the host of the heavens, those who bow down and swear to the LORD and yet swear by Milcom,
ZEPH|1|6|those who have turned back from following the LORD, who do not seek the LORD or inquire of him."
ZEPH|1|7|Be silent before the Lord GOD! For the day of the LORD is near; the LORD has prepared a sacrifice and consecrated his guests.
ZEPH|1|8|And on the day of the LORD's sacrifice- "I will punish the officials and the king's sons and all who array themselves in foreign attire.
ZEPH|1|9|On that day I will punish everyone who leaps over the threshold, and those who fill their master's house with violence and fraud.
ZEPH|1|10|"On that day," declares the LORD, "a cry will be heard from the Fish Gate, a wail from the Second Quarter, a loud crash from the hills.
ZEPH|1|11|Wail, O inhabitants of the Mortar! For all the traders are no more; all who weigh out silver are cut off.
ZEPH|1|12|At that time I will search Jerusalem with lamps, and I will punish the men who are complacent, those who say in their hearts, 'The LORD will not do good, nor will he do ill.'
ZEPH|1|13|Their goods shall be plundered, and their houses laid waste. Though they build houses, they shall not inhabit them; though they plant vineyards, they shall not drink wine from them."
ZEPH|1|14|The great day of the LORD is near, near and hastening fast; the sound of the day of the LORD is bitter; the mighty man cries aloud there.
ZEPH|1|15|A day of wrath is that day, a day of distress and anguish, a day of ruin and devastation, a day of darkness and gloom, a day of clouds and thick darkness,
ZEPH|1|16|a day of trumpet blast and battle cry against the fortified cities and against the lofty battlements.
ZEPH|1|17|I will bring distress on mankind, so that they shall walk like the blind, because they have sinned against the LORD; their blood shall be poured out like dust, and their flesh like dung.
ZEPH|1|18|Neither their silver nor their gold shall be able to deliver them on the day of the wrath of the LORD. In the fire of his jealousy, all the earth shall be consumed; for a full and sudden end he will make of all the inhabitants of the earth.
ZEPH|2|1|Gather together, yes, gather, O shameless nation,
ZEPH|2|2|before the decree takes effect- before the day passes away like chaff- before there comes upon you the burning anger of the LORD, before there comes upon you the day of the anger of the LORD.
ZEPH|2|3|Seek the LORD, all you humble of the land, who do his just commands; seek righteousness; seek humility; perhaps you may be hidden on the day of the anger of the LORD.
ZEPH|2|4|For Gaza shall be deserted, and Ashkelon shall become a desolation; Ashdod's people shall be driven out at noon, and Ekron shall be uprooted.
ZEPH|2|5|Woe to you inhabitants of the seacoast, you nation of the Cherethites! The word of the LORD is against you, O Canaan, land of the Philistines; and I will destroy you until no inhabitant is left.
ZEPH|2|6|And you, O seacoast, shall be pastures, with meadows for shepherds and folds for flocks.
ZEPH|2|7|The seacoast shall become the possession of the remnant of the house of Judah, on which they shall graze, and in the houses of Ashkelon they shall lie down at evening. For the LORD their God will be mindful of them and restore their fortunes.
ZEPH|2|8|"I have heard the taunts of Moab and the revilings of the Ammonites, how they have taunted my people and made boasts against their territory.
ZEPH|2|9|Therefore, as I live," declares the LORD of hosts, the God of Israel, "Moab shall become like Sodom, and the Ammonites like Gomorrah, a land possessed by nettles and salt pits, and a waste forever. The remnant of my people shall plunder them, and the survivors of my nation shall possess them."
ZEPH|2|10|This shall be their lot in return for their pride, because they taunted and boasted against the people of the LORD of hosts.
ZEPH|2|11|The LORD will be awesome against them; for he will famish all the gods of the earth, and to him shall bow down, each in its place, all the lands of the nations.
ZEPH|2|12|You also, O Cushites, shall be slain by my sword.
ZEPH|2|13|And he will stretch out his hand against the north and destroy Assyria, and he will make Nineveh a desolation, a dry waste like the desert.
ZEPH|2|14|Herds shall lie down in her midst, all kinds of beasts; even the owl and the hedgehog shall lodge in her capitals; a voice shall hoot in the window; devastation will be on the threshold; for her cedar work will be laid bare.
ZEPH|2|15|This is the exultant city that lived securely, that said in her heart, "I am, and there is no one else." What a desolation she has become, a lair for wild beasts! Everyone who passes by her hisses and shakes his fist.
ZEPH|3|1|Woe to her who is rebellious and defiled, the oppressing city!
ZEPH|3|2|She listens to no voice; she accepts no correction. She does not trust in the LORD; she does not draw near to her God.
ZEPH|3|3|Her officials within her are roaring lions; her judges are evening wolves that leave nothing till the morning.
ZEPH|3|4|Her prophets are fickle, treacherous men; her priests profane what is holy; they do violence to the law.
ZEPH|3|5|The LORD within her is righteous; he does no injustice; every morning he shows forth his justice; each dawn he does not fail; but the unjust knows no shame.
ZEPH|3|6|"I have cut off nations; their battlements are in ruins; I have laid waste their streets so that no one walks in them; their cities have been made desolate, without a man, without an inhabitant.
ZEPH|3|7|I said, 'Surely you will fear me; you will accept correction. Then your dwelling would not be cut off according to all that I have appointed against you.' But all the more they were eager to make all their deeds corrupt.
ZEPH|3|8|"Therefore wait for me," declares the LORD, "for the day when I rise up to seize the prey. For my decision is to gather nations, to assemble kingdoms, to pour out upon them my indignation, all my burning anger; for in the fire of my jealousy all the earth shall be consumed.
ZEPH|3|9|"For at that time I will change the speech of the peoples to a pure speech, that all of them may call upon the name of the LORD and serve him with one accord.
ZEPH|3|10|From beyond the rivers of Cush my worshipers, the daughter of my dispersed ones, shall bring my offering.
ZEPH|3|11|"On that day you shall not be put to shame because of the deeds by which you have rebelled against me; for then I will remove from your midst your proudly exultant ones, and you shall no longer be haughty in my holy mountain.
ZEPH|3|12|But I will leave in your midst a people humble and lowly. They shall seek refuge in the name of the LORD,
ZEPH|3|13|those who are left in Israel; they shall do no injustice and speak no lies, nor shall there be found in their mouth a deceitful tongue. For they shall graze and lie down, and none shall make them afraid."
ZEPH|3|14|Sing aloud, O daughter of Zion; shout, O Israel! Rejoice and exult with all your heart, O daughter of Jerusalem!
ZEPH|3|15|The LORD has taken away the judgments against you; he has cleared away your enemies. The King of Israel, the LORD, is in your midst; you shall never again fear evil.
ZEPH|3|16|On that day it shall be said to Jerusalem: "Fear not, O Zion; let not your hands grow weak.
ZEPH|3|17|The LORD your God is in your midst, a mighty one who will save; he will rejoice over you with gladness; he will quiet you by his love; he will exult over you with loud singing.
ZEPH|3|18|I will gather those of you who mourn for the festival, so that you will no longer suffer reproach.
ZEPH|3|19|Behold, at that time I will deal with all your oppressors. And I will save the lame and gather the outcast, and I will change their shame into praise and renown in all the earth.
ZEPH|3|20|At that time I will bring you in, at the time when I gather you together; for I will make you renowned and praised among all the peoples of the earth, when I restore your fortunes before your eyes," says the LORD.
