2SAM|1|1|Factum est autem, postquam mortuus est Saul, ut David re verteretur a caede Amalec et maneret in Siceleg dies duos.
2SAM|1|2|In die autem tertia apparuit homo veniens de castris Saul veste conscissa et pulvere aspersus caput; et, ut venit ad David, cecidit super faciem suam et adoravit.
2SAM|1|3|Dixitque ad eum David: " Unde venis? ". Qui ait ad eum: " De castris Israel fugi ".
2SAM|1|4|Et dixit ad eum David: " Quid enim factum est? Indica mihi ". Qui ait: " Fugit populus ex proelio, et multi corruentes e populo mortui sunt; sed et Saul et Ionathan filius eius interierunt ".
2SAM|1|5|Dixitque David ad adulescentem, qui nuntiabat ei: " Unde scis quia mortuus est Saul et Ionathan filius eius? ".
2SAM|1|6|Et ait adulescens, qui narrabat ei: " Casu veni in montem Gelboe, et Saul incumbebat super hastam suam. Porro currus et equites appropinquabant ei,
2SAM|1|7|et conversus post tergum suum vidensque me vocavit. Cui cum respondissem: Adsum,
2SAM|1|8|dixit mihi: "Quisnam es tu?". Et dixi ad eum: Amalecites ego sum.
2SAM|1|9|Et locutus est mihi: "Sta super me et interfice me, quoniam tenent me angustiae, et adhuc tota anima mea in me est".
2SAM|1|10|Stansque super eum occidi illum; sciebam enim quod vivere non poterat post ruinam. Et tuli diadema, quod erat in capite eius, et armillam de brachio illius et attuli ad te dominum meum huc ".
2SAM|1|11|Apprehendens autem David vestimenta sua scidit omnesque viri, qui erant cum eo;
2SAM|1|12|et planxerunt et fleverunt et ieiunaverunt usque ad vesperam super Saul et super Ionathan filium eius et super populum Domini et super domum Israel, quod corruissent gladio.
2SAM|1|13|Dixitque David ad iuvenem, qui nuntiaverat ei: " Unde es? ". Qui respondit: " Filius hominis advenae Amalecitae ego sum ".
2SAM|1|14|Et ait ad eum David: " Quare non timuisti mittere manum tuam, ut occideres christum Domini? ".
2SAM|1|15|Vocansque David unum de pueris ait: " Accedens irrue in eum ". Qui percussit illum, et mortuus est.
2SAM|1|16|Et ait ad eum David: " Sanguis tuus super caput tuum; os enim tuum locutum est adversum te dicens: "Ego interfeci christum Domini" ".
2SAM|1|17|Planxit autem David planctum huiuscemodi super Saul et super Ionathan filium eius;
2SAM|1|18|et praecepit, ut docerent filios Iudae canticum Arcus, sicut scriptum est in libro Iusti, et ait:
2SAM|1|19|" Incliti, o Israel, super montes tuos interfecti,quomodo ceciderunt fortes!
2SAM|1|20|Nolite annuntiare in Gethneque annuntietis in compitis Ascalonis,ne forte laetentur filiae Philisthim,ne exsultent filiae incircumcisorum.
2SAM|1|21|Montes Gelboe, nec ros nec pluviae veniant super vos,neque sint agri oblationum!Quia ibi abiectus est clipeus fortium,clipeus Saul, quasi non esset unctus oleo.
2SAM|1|22|A sanguine interfectorum, ab adipe fortiumarcus Ionathan numquam rediit retrorsum,et gladius Saul non est reversus inanis.
2SAM|1|23|Saul et Ionathan amabiles et decori in vita sua,in morte quoque non sunt divisi,aquilis velociores, leonibus fortiores.
2SAM|1|24|Filiae Israel, super Saul flete,qui vestiebat vos coccino in deliciis, qui praebebat ornamenta aurea cultui vestro.
2SAM|1|25|Quomodo ceciderunt fortes in proelio!Ionathan in excelsis tuis occisus est.
2SAM|1|26|Doleo super te, frater mi Ionathan,suavis nimis mihi;mirabilis amor tuus mihisuper amorem mulierum.
2SAM|1|27|Quomodo ceciderunt fortes,et perierunt arma bellica! ".
2SAM|2|1|Igitur post haec consuluit David Dominum dicens: " Num ascendam in unam de civitatibus Iudae? ". Et ait Dominus ad eum: " Ascende ". Dixitque David: " Quo ascendam? ". Et respondit ei: " In Hebron ".
2SAM|2|2|Ascendit ergo David et duae uxores eius, Achinoam Iezrahelites et Abigail uxor Nabal de Carmel;
2SAM|2|3|sed et viros, qui erant cum eo, duxit David singulos cum domo sua, et manserunt in oppidis Hebron.
2SAM|2|4|Veneruntque viri Iudae et unxerunt ibi David, ut regnaret super domum Iudae.Et nuntiatum est David quod viri Iabes Galaad sepelissent Saul.
2SAM|2|5|Misit ergo David nuntios ad viros Iabes Galaad dixitque ad eos: " Benedicti vos Domino, qui fecistis misericordiam hanc cum domino vestro Saul et sepelistis eum.
2SAM|2|6|Et nunc faciat quidem vobis Dominus misericordiam et veritatem; sed et ego reddam vobis similiter bonum, eo quod feceritis istud.
2SAM|2|7|Nunc autem confortentur manus vestrae, et estote fortes; licet enim mortuus sit dominus vester Saul, tamen me unxit domus Iudae in regem sibi.
2SAM|2|8|Abner autem filius Ner princeps exercitus Saul tulit Isbaal filium Saul et duxit eum in Mahanaim
2SAM|2|9|regemque constituit super Galaad et super Aser et super Iezrahel et super Ephraim et super Beniamin et super Israel universum.
2SAM|2|10|Quadraginta annorum erat Isbaal filius Saul, cum regnare coepisset super Israel, et duobus annis regnavit; sola autem domus Iudae sequebatur David.
2SAM|2|11|Et fuit numerus dierum, quos commoratus est David imperans in Hebron super domum Iudae, septem annorum et sex mensium.
2SAM|2|12|Egressusque est Abner filius Ner et pueri Isbaal filii Saul de Mahanaim in Gabaon.
2SAM|2|13|Porro Ioab filius Sarviae et pueri David egressi sunt et occurrerunt eis iuxta piscinam Gabaon; et, cum in unum convenissent e regione, constiterunt hi ex una parte piscinae et illi ex altera.
2SAM|2|14|Dixitque Abner ad Ioab: " Surgant pueri et ludant coram nobis ". Et respondit Ioab: " Surgant ".
2SAM|2|15|Surrexerunt ergo et transierunt numero duodecim de Beniamin ex parte Isbaal filii Saul, et duodecim de pueris David.
2SAM|2|16|Apprehensoque unusquisque capite comparis sui, defixit gladium in latus contrarii, et ceciderunt simul; vocatumque est nomen loci illius ager Laterum in Gabaon.
2SAM|2|17|Et ortum est bellum durum valde in die illa, fugatusque est Abner et viri Israel a pueris David.
2SAM|2|18|Erant autem ibi tres filii Sarviae: Ioab et Abisai et Asael. Porro Asael cursor velocissimus fuit quasi unus ex capreis, quae morantur in campis.
2SAM|2|19|Persequebatur autem Asael Abner et non declinavit ad dextram sive ad sinistram omittens persequi Abner.
2SAM|2|20|Respexit itaque Abner post tergum suum et ait: " Tune es Asael? ". Qui respondit: " Ego sum ".
2SAM|2|21|Dixitque ei Abner: " Vade ad dextram sive ad sinistram et apprehende unum de adulescentibus et tolle tibi spolia eius ". Noluit autem Asael omittere quin urgeret eum.
2SAM|2|22|Rursumque locutus est Abner ad Asael: " Recede, noli me sequi, ne compellar confodere te in terram et levare non potero faciem meam ad Ioab fratrem tuum ".
2SAM|2|23|Qui audire contempsit et noluit declinare. Percussit ergo eum Abner, aversa hasta in inguine, et exiit hasta retrorsum, et mortuus est ibi. Omnesque qui transibant per locum, in quo ceciderat Asael et mortuus erat, subsistebant.
2SAM|2|24|Persequentibus autem Ioab et Abisai fugientem Abner, sol occubuit; et venerunt usque ad collem Amma, qui est ex adverso Gaiah in via deserti in Gabaon.
2SAM|2|25|Congregatique sunt filii Beniamin ad Abner et conglobati in unum cuneum steterunt in summitate tumuli unius.
2SAM|2|26|Et exclamavit Abner ad Ioab et ait: " Num usque ad internecionem tuus mucro desaeviet? An ignoras quod periculosa sit desperatio? Usquequo non dicis populo, ut omittat persequi fratres suos? ".
2SAM|2|27|Et ait Ioab: " Vivit Deus, nisi locutus fuisses, usque mane non recessisset populus persequens unusquisque fratrem suum ".
2SAM|2|28|Insonuit ergo Ioab bucina, et stetit omnis exercitus; nec persecuti sunt ultra Israel neque certaverunt amplius.
2SAM|2|29|Abner autem et viri eius abierunt per Arabam tota nocte illa et transierunt Iordanem et, lustrato toto saltu Bethron, venerunt Mahanaim.
2SAM|2|30|Porro Ioab reversus, omisso Abner, congregavit omnem populum; et defuerunt de pueris David decem et novem viri, excepto Asaele;
2SAM|2|31|servi autem David percusserunt de Beniamin et ex viris, qui erant cum Abner, trecentos sexaginta, qui et mortui sunt.
2SAM|2|32|Tuleruntque Asael et sepelierunt eum in sepulcro patris sui in Bethlehem. Et ambulaverunt tota nocte Ioab et viri, qui erant cum eo, et in ipso crepusculo pervenerunt in Hebron.
2SAM|3|1|Facta est ergo longa concertatio inter domum Saul et inter do mum David: David semper invalescens, domus autem Saul decrescens cotidie.
2SAM|3|2|Nati quoque sunt filii David in Hebron. Fuitque primogenitus eius Amnon de Achinoam Iezrahelitide,
2SAM|3|3|et post eum Cheleab de Abigail uxore Nabal de Carmel, porro tertius Absalom filius Maacha filiae Tholmai regis Gesur,
2SAM|3|4|quartus autem Adonias filius Haggith et quintus Saphatia filius Abital,
2SAM|3|5|sextus quoque Iethraam de Egla uxore David. Hi nati sunt David in Hebron.
2SAM|3|6|Cum ergo esset proelium inter domum Saul et domum David, Abner filius Ner regebat domum Saul.
2SAM|3|7|Fuerat autem Sauli concubina nomine Respha filia Aia. Dixitque Isbaal ad Abner:
2SAM|3|8|" Quare ingressus es ad concubinam patris mei? ". Qui iratus nimis propter verba Isbaal ait: " Numquid caput canis ego sum de Iuda? Hodie facio misericordiam super domum Saul patris tui et super fratres et proximos eius et non tradidi te in manu David. Et tu requisisti in me quod argueres pro muliere hodie.
2SAM|3|9|Haec faciat Deus Abner et haec addat ei, nisi, quomodo iuravit Dominus David, sic faciam cum eo,
2SAM|3|10|ut transferatur regnum de domo Saul, et confirmetur thronus David super Israel et super Iudam a Dan usque Bersabee ".
2SAM|3|11|Et non potuit respondere ei quidquam, quia metuebat illum.
2SAM|3|12|Misit ergo Abner nuntios ad David pro se dicentes: " Cuius est terra?, et ut loquerentur: " Fac mecum amicitias, et erit manus mea tecum, et reducam ad te universum Israel ".
2SAM|3|13|Qui ait: " Optime, ego faciam tecum amicitias, sed unam rem peto a te dicens: Non videbis faciem meam, nisi prius adduxeris Michol filiam Saul; et sic venies et videbis me ".
2SAM|3|14|Misit autem David nuntios ad Isbaal filium Saul dicens: "Redde uxorem meam Michol, quam despondi mihi centum praeputiis Philisthim ".
2SAM|3|15|Misit ergo Isbaal et tulit eam a viro suo Phaltiel filio Lais.
2SAM|3|16|Sequebaturque eam vir suus plorans usque Bahurim; et dixit ad eum Abner: " Vade, revertere ". Qui reversus est.
2SAM|3|17|Sermonem quoque intulit Abner ad seniores Israel dicens: " Tam heri quam nudiustertius quaerebatis David, ut regnaret super vos;
2SAM|3|18|nunc ergo facite, quoniam Dominus locutus est ad David dicens: "In manu servi mei David salvabo populum meum Israel de manu Philisthim et omnium inimicorum eius" ".
2SAM|3|19|Locutus est autem Abner etiam ad Beniamin; et abiit, ut loqueretur ad David in Hebron omnia, quae placuerant Israel et universo Beniamin.
2SAM|3|20|Venitque ad David in Hebron cum viginti viris, et fecit David Abner et viris eius, qui venerant cum eo, convivium.
2SAM|3|21|Et dixit Abner ad David: " Surgam, ut congregem ad te dominum meum regem omnem Israel, et ineant tecum foedus, et imperes omnibus, sicut desiderat anima tua ".Cum ergo deduxisset David Abner, et ille isset in pace,
2SAM|3|22|pueri David et Ioab venerunt ab expeditione cum praeda magna. Abner autem non erat cum David in Hebron, quia iam dimiserat eum, et profectus fuerat in pace,
2SAM|3|23|et Ioab et omnis exercitus, qui erat cum eo, postea venerant. Nuntiatum est itaque Ioab a narrantibus: " Venit Abner filius Ner ad regem, et dimisit eum, et abiit in pace ".
2SAM|3|24|Et ingressus est Ioab ad regem et ait: " Quid fecisti? Ecce venit Abner ad te; quare dimisisti eum, et abiit et recessit?
2SAM|3|25|Ignoras Abner filium Ner? Certe ad hoc venit, ut deciperet te et sciret exitum tuum et introitum tuum et nosset omnia quae agis ".
2SAM|3|26|Egressus itaque Ioab a David misit nuntios post Abner, et reduxerunt eum a cisterna Sira, ignorante David.
2SAM|3|27|Cumque redisset Abner in Hebron, seorsum abduxit eum Ioab ad medium portae, ut loqueretur ei quiete, et percussit illum ibi in inguine, et mortuus est in ultionem sanguinis Asael fratris eius.
2SAM|3|28|Quod cum audisset David rem iam gestam, ait: " Mundus ego sum et regnum meum apud Dominum usque in sempiternum a sanguine Abner filii Ner;
2SAM|3|29|et veniat super caput Ioab et super omnem domum patris eius, nec deficiat de domo Ioab fluxum morbidum sustinens, leprosus et tenens fusum et cadens gladio et indigens pane ".
2SAM|3|30|Igitur Ioab et Abisai frater eius interfecerunt Abner, eo quod occidisset Asael fratrem eorum in Gabaon in proelio.
2SAM|3|31|Dixit autem David ad Ioab et ad omnem populum, qui erat cum eo: " Scindite vestimenta vestra et accingimini saccis et plangite ante exequias Abner ". Porro rex David sequebatur feretrum.
2SAM|3|32|Cumque sepelissent Abner in Hebron, levavit rex David vocem suam et flevit super tumulum Abner; flevit autem et omnis populus.
2SAM|3|33|Plangensque rex et lugens Abner ait: Numquid, ut mori solent insensati,mori debuit Abner?
2SAM|3|34|Manus tuae ligatae non erant,et pedes tui non erant compedibus aggravati;sed, sicut solent cadere coram filiis iniquitatis, corruisti ".Congeminansque omnis populus flevit super eum.
2SAM|3|35|Cumque venisset universa multitudo reficere David pane clara adhuc die, iuravit David dicens: " Haec faciat mihi Deus et haec addat, si ante occasum solis gustavero panem vel aliud quidquam ".
2SAM|3|36|Omnisque populus audivit; et placuit eis, sicut cuncta, quae fecit rex, bona erant in conspectu totius populi.
2SAM|3|37|Et cognovit omne vulgus et universus Israel in die illa quoniam non actum fuisset a rege, ut occideretur Abner filius Ner.
2SAM|3|38|Dixit quoque rex ad servos suos: " Num ignoratis quoniam princeps et maximus cecidit hodie in Israel?
2SAM|3|39|Ego vero adhuc debilis sum, quamvis sim unctus rex; viri autem isti filii Sarviae duriores sunt quam ego. Retribuat Dominus facienti malum iuxta malitiam suam ".
2SAM|4|1|Audivit autem Isbaal filius Saul quod cecidisset Abner in He bron, et dissolutae sunt manus eius, omnisque Israel perturbatus est.
2SAM|4|2|Duo autem viri duces turmarum erant filio Saul, nomen uni Baana et nomen alteri Rechab filii Remmon Berothitae de filiis Beniamin; siquidem et Beroth reputata est in Beniamin.
2SAM|4|3|Fugerant enim Berothitae in Getthaim, factique sunt ibi advenae usque in tempus hoc.
2SAM|4|4|Erat autem Ionathan filio Saul filius debilis pedibus. Quinquennis enim fuit, quando venit nuntius de Saul et Ionathan ex Iezrahel. Tollens itaque eum nutrix sua fugit; cumque festinaret, ut fugeret, cecidit et claudus effectus est habuitque vocabulum Meribbaal.
2SAM|4|5|Venientes igitur filii Remmon Berothitae, Rechab et Baana, ingressi sunt, fervente die, domum Isbaal, qui dormiebat super stratum suum meridie; et ostiaria domus purgans triticum obdormivit.
2SAM|4|6|Ingressi sunt ergo usque interiora domus et percusserunt eum in inguine Rechab et Baana frater eius et fugerunt.
2SAM|4|7|Cum autem ingressi fuissent domum, ille dormiebat super lectum suum in conclavi, et percutientes interfecerunt eum; sublatoque capite eius, abierunt per viam Arabae tota nocte.
2SAM|4|8|Et attulerunt caput Isbaal ad David in Hebron dixeruntque ad regem: " Ecce caput Isbaal filii Saul inimici tui, qui quaerebat animam tuam; et dedit Dominus domino meo regi ultiones hodie de Saul et de semine eius ".
2SAM|4|9|Respondens autem David Rechab et Baana fratri eius filiis Remmon Berothitae dixit ad eos: " Vivit Dominus, qui eruit animam meam de omni angustia,
2SAM|4|10|quoniam eum, qui annuntiaverat mihi et dixerat: "Mortuus est Saul", qui putabat se prospera nuntiare, tenui et occidi in Siceleg, cui oportebat me dare mercedem pro nuntio;
2SAM|4|11|quanto magis nunc, cum homines impii interfecerunt virum innoxium in domo sua super lectum suum, non quaeram sanguinem eius de manu vestra et auferam vos de terra? ".
2SAM|4|12|Praecepit itaque David pueris, et interfecerunt eos; praecidentesque manus et pedes eorum suspenderunt eos super piscinam in Hebron. Caput autem Isbaal tulerunt et sepelierunt in sepulcro Abner in Hebron.
2SAM|5|1|Et venerunt universae tribus Is rael ad David in Hebron dicen tes: " Ecce nos os tuum et caro tua sumus.
2SAM|5|2|Sed et heri et nudiustertius, cum esset Saul rex super nos, tu eras educens et reducens Israel. Dixit autem Dominus ad te: "Tu pasces populum meum Israel et tu eris dux super Israel" ".
2SAM|5|3|Venerunt quoque omnes senes Israel ad regem in Hebron, et percussit cum eis rex David foedus in Hebron coram Domino; unxeruntque David in regem super Israel.
2SAM|5|4|Triginta annorum erat David, cum regnare coepisset, et quadraginta annis regnavit:
2SAM|5|5|in Hebron regnavit super Iudam septem annis et sex mensibus; in Ierusalem autem regnavit triginta tribus annis super omnem Israel et Iudam.
2SAM|5|6|Et abiit rex et omnes viri, qui erant cum eo, in Ierusalem ad Iebusaeum habitatorem terrae. Qui dixit ad David: "Non ingredieris huc, sed depellent te caeci et claudi ", significantes: " Non ingredietur David huc.
2SAM|5|7|Cepit autem David arcem Sion: haec est civitas David.
2SAM|5|8|Dixerat enim David in die illa: " Omnis, qui percutiet Iebusaeum, attingat per cuniculum fontis claudos et caecos exosos animae David ". Idcirco dicitur in proverbio: " Caecus et claudus non intrabunt in domum.
2SAM|5|9|Habitavit autem David in arce et vocavit eam Civitatem David; et aedificavit per gyrum a Mello et intrinsecus.
2SAM|5|10|Et ibat proficiens atque succrescens, et Dominus, Deus exercituum, erat cum eo.
2SAM|5|11|Misit quoque Hiram rex Tyri nuntios ad David et ligna cedrina et artifices lignorum artificesque lapidum pro parietibus; et aedificaverunt domum David.
2SAM|5|12|Et cognovit David quoniam confirmasset eum Dominus regem super Israel et quoniam exaltasset regnum eius super populum suum Israel.
2SAM|5|13|Accepitque David adhuc concubinas et uxores de Ierusalem, postquam venerat de Hebron; natique sunt David et alii filii et filiae.
2SAM|5|14|Et haec nomina eorum, qui nati sunt ei in Ierusalem: Samua et Sobab et Nathan et Salomon
2SAM|5|15|et Iebahar et Elisua et Napheg
2SAM|5|16|et Iaphia et Elisama et Eliada et Eliphalet.
2SAM|5|17|Audierunt vero Philisthim quod unxissent David regem super Israel et ascenderunt universi, ut quaererent David. Quod cum audisset David, descendit in praesidium;
2SAM|5|18|Philisthim autem venientes diffusi sunt in valle Raphaim.
2SAM|5|19|Et consuluit David Dominum dicens: " Si ascendam ad Philisthim? Et si dabis eos in manu mea? ". Et dixit Dominus ad David: "Ascende, quia tradens dabo Philisthim in manu tua ".
2SAM|5|20|Venit ergo David in Baalpharasim (id est Dominus diruptionum); et percussit eos ibi et dixit: "Divisit Dominus inimicos meos coram me, sicut dividuntur aquae ". Propterea vocatum est nomen loci illius Baalpharasim.
2SAM|5|21|Et reliquerunt ibi sculptilia sua, quae tulit David et viri eius.
2SAM|5|22|Et addiderunt adhuc Philisthim ut ascenderent et diffusi sunt in valle Raphaim.
2SAM|5|23|Consuluit autem David Dominum, qui respondit: " Non ascendas, sed gyra post tergum eorum et venies ad eos ex adverso arborum celthium
2SAM|5|24|et, cum audieris sonitum gradientis in cacumine arborum celthium, tunc inibis proelium, quia tunc egredietur Dominus ante faciem tuam, ut percutiat castra Philisthim ".
2SAM|5|25|Fecit itaque David, sicut praeceperat ei Dominus; et percussit Philisthim de Gabaon usque dum venias Gazer.
2SAM|6|1|Congregavit autem rursum Da vid omnes electos ex Israel tri ginta milia.
2SAM|6|2|Surrexitque David et abiit, et universus populus, qui erat cum eo, in Baala Iudae, ut adducerent inde arcam Dei, super quam invocatum est nomen Domini exercituum sedentis in cherubim super eam.
2SAM|6|3|Et imposuerunt arcam Dei super plaustrum novum tuleruntque eam de domo Abinadab, qui erat in colle. Oza autem et Ahio filii Abinadab minabant plaustrum:
2SAM|6|4|Oza ambulabat iuxta arcam, et Ahio praecedebat eam.
2SAM|6|5|David autem et omnis Israel ludebant coram Domino omni virtute in canticis et citharis et lyris et tympanis et sistris et cymbalis.
2SAM|6|6|Postquam autem venerunt ad aream Nachon, extendit manum Oza ad arcam Dei et tenuit eam, quoniam boves lascivientes proruperunt.
2SAM|6|7|Iratusque est indignatione Dominus contra Ozam et percussit eum super temeritate; qui mortuus est ibi iuxta arcam Dei.
2SAM|6|8|Contristatus autem est David, eo quod diruptionem dirupisset Dominus in Ozam; et vocatum est nomen loci illius Pharesoza (id est Diruptio Ozae) usque in diem hanc.
2SAM|6|9|Et extimuit David Dominum in die illa dicens: " Quomodo ingredietur ad me arca Domini? ".
2SAM|6|10|Et noluit divertere ad se arcam Domini in civitate David, sed divertit eam in domum Obededom Getthaei.
2SAM|6|11|Et habitavit arca Domini in domo Obededom Getthaei tribus mensibus, et benedixit Dominus Obededom et omnem domum eius.
2SAM|6|12|Nuntiatumque est regi David: " Benedixit Dominus Obededom et omnia eius propter arcam Dei ". Abiit ergo David et adduxit arcam Dei de domo Obededom in civitatem David cum gaudio.
2SAM|6|13|Cumque progressi essent, qui portabant arcam Domini, sex passus, immolavit bovem et vitulum saginatum,
2SAM|6|14|et David saltabat totis viribus ante Dominum. Porro David erat accinctus ephod lineo.
2SAM|6|15|Et David et omnis domus Israel ducebant arcam Domini in iubilo et in clangore bucinae.
2SAM|6|16|Cumque intrasset arca Domini in civitatem David, Michol filia Saul prospiciens per fenestram vidit regem David subsilientem atque saltantem coram Domino et despexit eum in corde suo.
2SAM|6|17|Et introduxerunt arcam Domini et posuerunt eam in loco suo in medio tabernaculi, quod tetenderat ei David; et obtulit David coram Domino holocausta et pacifica.
2SAM|6|18|Cumque complesset offerens holocaustum et pacifica, benedixit populo in nomine Domini exercituum.
2SAM|6|19|Et partitus est multitudini universae Israel tam viro quam mulieri singulis collyridam panis unam et laganum palmarum unum et palatham unam. Et abiit omnis populus unusquisque in domum suam.
2SAM|6|20|Reversusque est et David, ut benediceret domui suae, et egressa Michol filia Saul in occursum David ait: " Quam gloriosus fuit hodie rex Israel discooperiens se ante ancillas servorum suorum, quasi si nudetur unus de scurris! ".
2SAM|6|21|Dixitque David ad Michol: " Ante Dominum salto. Benedictus Dominus, qui elegit me potius quam patrem tuum et quam omnem domum eius, ut constitueret me ducem super populum Domini, super Israel!
2SAM|6|22|Ludam in conspectu Domini et vilior fiam plus quam factus sum et ero deiectus in oculis meis, sed apud ancillas, de quibus locuta es, gloriosior apparebo ".
2SAM|6|23|Igitur Michol filiae Saul non est natus filius usque ad diem mortis suae.
2SAM|7|1|Factum est autem cum sedisset rex in domo sua, et Dominus de disset ei requiem undique ab universis inimicis suis,
2SAM|7|2|dixit ad Nathan prophetam: " Videsne quod ego habitem in domo cedrina, et arca Dei posita sit in medio pellium? ".
2SAM|7|3|Dixitque Nathan ad regem: " Omne, quod est in corde tuo, vade, fac, quia Dominus tecum est ".
2SAM|7|4|Factum est autem in nocte illa, et ecce sermo Domini ad Nathan dicens:
2SAM|7|5|" Vade et loquere ad servum meum David: Haec dicit Dominus: Numquid tu aedificabis mihi domum ad habitandum?
2SAM|7|6|Numquam enim habitavi in domo ex die, qua eduxi filios Israel de terra Aegypti, usque in diem hanc, sed ambulabam in tabernaculo et in tentorio.
2SAM|7|7|Per cuncta loca, quae transivi cum omnibus filiis Israel, numquid loquens locutus sum ad unum de iudicibus Israel, cui praecepi, ut pasceret populum meum Israel, dicens: Quare non aedificastis mihi domum cedrinam?
2SAM|7|8|Et nunc haec dices servo meo David: Haec dicit Dominus exercituum: Ego tuli te de pascuis sequentem greges, ut esses dux super populum meum Israel,
2SAM|7|9|et fui tecum in omnibus, ubicumque ambulasti, et interfeci universos inimicos tuos a facie tua; fecique tibi nomen grande iuxta nomen magnorum, qui sunt in terra.
2SAM|7|10|Et ponam locum populo meo Israel et plantabo eum, et habitabit in eo et non turbabitur amplius; nec addent filii iniquitatis ut affligant eum sicut prius
2SAM|7|11|et ex die, qua constitui iudices super populum meum Israel, et requiem dabo tibi ab omnibus inimicis tuis. Praedicitque tibi Dominus quod domum faciat tibi Dominus.
2SAM|7|12|Cumque completi fuerint dies tui, et dormieris cum patribus tuis, suscitabo semen tuum post te, quod egredietur de visceribus tuis; et firmabo regnum eius.
2SAM|7|13|Ipse aedificabit domum nomini meo, et stabiliam thronum regni eius usque in sempiternum.
2SAM|7|14|Ego ero ei in patrem, et ipse erit mihi in filium; qui si inique aliquid gesserit, arguam eum in virga virorum et in plagis filiorum hominum.
2SAM|7|15|Misericordiam autem meam non auferam ab eo, sicut abstuli a Saul, quem amovi a facie tua;
2SAM|7|16|et stabilis erit domus tua et regnum tuum usque in aeternum ante faciem meam, et thronus tuus erit firmus iugiter ".
2SAM|7|17|Secundum omnia verba haec et iuxta universam visionem istam sic locutus est Nathan ad David.
2SAM|7|18|Ingressus est autem rex David et sedit coram Domino et dixit: " Quis ego sum, Domine Deus, et quae domus mea, quia adduxisti me hucusque?
2SAM|7|19|Sed et hoc parum visum est in conspectu tuo, Domine Deus, et locutus es etiam de domo servi tui in longinquum, et ista est lex hominis, Domine Deus!
2SAM|7|20|Quid ergo addere poterit adhuc David, ut loquatur ad te? Tu enim scis servum tuum, Domine Deus.
2SAM|7|21|Propter verbum tuum et secundum cor tuum fecisti omnia magnalia haec, ita ut nota faceres servo tuo.
2SAM|7|22|Idcirco magnus es, Domine Deus, quia non est similis tui; neque est Deus extra te, iuxta omnia, quae audivimus auribus nostris.
2SAM|7|23|Quae est autem ut populus tuus Israel una gens in terra, propter quam ivit Deus, ut redimeret eam sibi in populum et poneret sibi nomen faceretque eis magnalia et horribilia, ut eiceres a facie populi tui, quem redemisti tibi ex Aegypto, gentes et deos eorum?
2SAM|7|24|Et firmasti tibi populum tuum Israel in populum sempiternum; et tu, Domine, factus es eis in Deum.
2SAM|7|25|Nunc ergo, Domine Deus, verbum, quod locutus es super servum tuum et super domum eius, confirma in sempiternum et fac, sicut locutus es!
2SAM|7|26|Et magnificetur nomen tuum usque in sempiternum, atque dicatur: Dominus exercituum est Deus super Israel". Et domus servi tui David erit stabilita coram te,
2SAM|7|27|quia tu, Domine exercituum, Deus Israel, revelasti aurem servi tui dicens: "Domum aedificabo tibi". Propterea invenit servus tuus cor suum, ut oraret te oratione hac.
2SAM|7|28|Nunc ergo, Domine Deus, tu es Deus, et verba tua erunt vera; cum ergo locutus sis ad servum tuum bona haec,
2SAM|7|29|dignare igitur benedicere domui servi tui, ut sit in sempiternum coram te, quia tu, Domine Deus, locutus es, et benedictione tua benedicetur domus servi tui in sempiternum ".
2SAM|8|1|Factum est autem post haec, percussit David Philisthim et humiliavit eos; et tulit David Geth et urbes eius de manu Philisthim.
2SAM|8|2|Et percussit Moab et mensus est eos funiculo sternens eos in terra; mensus est autem duos funiculos ad occidendum et unum funiculum plenum ad vivificandum; factusque est Moab David serviens sub tributo.
2SAM|8|3|Et percussit David Adadezer filium Rohob regem Soba, quando profectus est, ut dominaretur super flumen Euphraten.
2SAM|8|4|Et captis David ex parte eius mille septingentis equitibus et viginti milibus peditum, subnervavit omnes iugales curruum; dereliquit autem ex eis centum currus.
2SAM|8|5|Venit quoque Syria Damasci, ut praesidium ferret Adadezer regi Soba, et percussit David de Syria viginti duo milia virorum;
2SAM|8|6|et posuit David praesidium in Syria Damasci; factaque est Syria David serviens sub tributo. Et auxiliatus est Dominus David in omnibus, ad quaecumque profectus est.
2SAM|8|7|Et tulit David arma aurea, quae habebant servi Adadezer, et detulit ea in Ierusalem;
2SAM|8|8|et de Tebah et de Berothai civitatibus Adadezer tulit rex David aes multum nimis.
2SAM|8|9|Audivit autem Thou rex Emath quod percussisset David omne robur Adadezer
2SAM|8|10|et misit Thou Adoram filium suum ad regem David, ut salutaret eum congratulans et gratias ageret eo quod pugnasset cum Adadezer et percussisset eum; hostis quippe erat Thou Adadezer. Attulit autem Adoram et vasa argentea et vasa aurea et vasa aerea,
2SAM|8|11|quae et ipsa sanctificavit rex David Domino cum argento et auro, quae sanctificaverat de universis gentibus, quas subegerat:
2SAM|8|12|de Syria et Moab et filiis Ammon et Philisthim et Amalec et de manibus Adadezer filii Rohob regis Soba.
2SAM|8|13|Fecit quoque sibi David nomen cum reverteretur, percussa Idumaea in valle Salis, caesis decem et octo milibus.
2SAM|8|14|Et posuit in Idumaea praesidia; et facta est universa Idumaea serviens David. Et auxiliatus est Dominus David in omnibus, ad quaecumque profectus est.
2SAM|8|15|Et regnavit David super omnem Israel; faciebat quoque David iudicium et iustitiam omni populo suo.
2SAM|8|16|Ioab autem filius Sarviae erat super exercitum; porro Iosaphat filius Ahilud erat a commentariis,
2SAM|8|17|et Sadoc filius Achitob et Abiathar filius Achimelech sacerdotes, et Saraias scriba.
2SAM|8|18|Banaias autem filius Ioiadae super Cherethi et Phelethi; filii autem David sacerdotes erant.
2SAM|9|1|Et dixit David: " Putasne est aliquis, qui remanserit adhuc de domo Saul, ut faciam cum eo misericordiam propter Ionathan? ".
2SAM|9|2|Erat autem de domo Saul servus nomine Siba; quem cum vocasset rex ad se, dixit ei: " Tune es Siba? ". Et ille respondit: " Ego sum, servus tuus ".
2SAM|9|3|Et ait rex: " Num superest aliquis de domo Saul, ut faciam cum eo misericordiam Dei? ". Dixitque Siba regi: " Superest filius Ionathan, debilis pedibus ".
2SAM|9|4|" Ubi, inquit, est? ". Et Siba ad regem: " Ecce, ait, in domo est Machir filii Ammiel in Lodabar ".
2SAM|9|5|Misit ergo rex David et tulit eum de domo Machir filii Ammiel de Lodabar.
2SAM|9|6|Cum autem venisset Meribbaal filius Ionathan filii Saul ad David, corruit in faciem suam et adoravit. Dixitque David: " Meribbaal ". Qui respondit: " Adsum servus tuus ".
2SAM|9|7|Et ait ei David: "Ne timeas, quia faciens faciam in te misericordiam propter Ionathan patrem tuum; et restituam tibi omnes agros Saul patris tui, et tu comedes panem in mensa mea semper ".
2SAM|9|8|Qui adorans eum dixit: " Quis ego sum servus tuus, quoniam respexisti super canem mortuum similem mei? ".
2SAM|9|9|Vocavit itaque rex Sibam puerum Saul et dixit ei: " Omnia, quaecumque fuerunt Saul et universae domui eius, do filio domini tui.
2SAM|9|10|Operare igitur ei terram, tu et filii tui et servi tui, et, quod inferes, sit cibus domui domini tui, quo alantur; Meribbaal autem filius domini tui comedet semper panem super mensam meam ". Erant autem Sibae quindecim filii et viginti servi.
2SAM|9|11|Dixitque Siba ad regem: " Sicut iussisti, domine mi rex, servo tuo, sic faciet servus tuus ". Meribbaal autem comedebat super mensam eius quasi unus de filiis regis.
2SAM|9|12|Habebat autem Meribbaal filium parvulum nomine Micha; omnes vero, qui habitabant in domo Sibae, serviebant Meribbaal.
2SAM|9|13|Porro Meribbaal habitabat in Ierusalem, quia de mensa regis iugiter vescebatur; et erat claudus utroque pede.
2SAM|10|1|Factum est autem post haec, ut moreretur rex filiorum Ammon, et regnaret Hanon filius eius pro eo.
2SAM|10|2|Dixitque David: " Faciam misericordiam cum Hanon filio Naas, sicut fecit pater eius mecum misericordiam ". Misit ergo David consolans eum per servos suos super patris interitu. Cum autem venissent servi David in terram filiorum Ammon,
2SAM|10|3|dixerunt principes filiorum Ammon ad Hanon dominum suum: " Putas quod propter honorem patris tui David miserit ad te consolatores; et non ideo, ut investigaret et exploraret civitatem et everteret eam, misit David servos suos ad te? ".
2SAM|10|4|Tulit itaque Hanon servos David rasitque dimidiam partem barbae eorum et praecidit vestes eorum medias usque ad nates et dimisit eos.
2SAM|10|5|Quod cum nuntiatum esset David, misit in occursum eorum - erant enim viri confusi turpiter valde - et mandavit eis David: " Manete Iericho, donec crescat barba vestra, et tunc revertimini ".
2SAM|10|6|Videntes autem filii Ammon quod exosos se fecissent David, miserunt et conduxerunt mercede a Syria Bethrohob et a Syria Soba viginti milia peditum et a rege Maacha mille viros et a viris Tob duodecim milia virorum.
2SAM|10|7|Quod cum audisset David, misit Ioab et omnem exercitum, viros fortissimos.
2SAM|10|8|Egressi sunt ergo filii Ammon et direxerunt aciem ante ipsum introitum portae; Syri autem Soba et Rohob et viri Tob et Maacha seorsum erant in campo.
2SAM|10|9|Videns igitur Ioab quod praeparatum esset adversum se proelium et ex adverso et post tergum, elegit ex omnibus electis Israel et instruxit aciem contra Syros;
2SAM|10|10|reliquam autem partem populi tradidit Abisai fratri suo, qui direxit aciem adversus filios Ammon.
2SAM|10|11|Et ait Ioab: " Si praevaluerint adversum me Syri, eris mihi in adiutorium; si autem filii Ammon praevaluerint adversum te, auxiliabor tibi.
2SAM|10|12|Esto vir fortis, et fortiter agamus pro populo nostro et civitatibus Dei nostri; Dominus autem faciet, quod bonum est in conspectu suo ".
2SAM|10|13|Iniit itaque Ioab et populus, qui erat cum eo, certamen contra Syros, qui fugerunt a facie eius.
2SAM|10|14|Filii autem Ammon videntes quod fugissent Syri, fugerunt et ipsi a facie Abisai et ingressi sunt civitatem. Reversusque est Ioab a filiis Ammon et venit Ierusalem.
2SAM|10|15|Videntes igitur Syri quoniam corruissent coram Israel, congregati sunt pariter.
2SAM|10|16|Misitque Adadezer et eduxit Syros, qui erant trans fluvium, et venerunt in Elam; Sobach autem magister militiae Adadezer erat princeps eorum.
2SAM|10|17|Quod cum nuntiatum esset David, contraxit omnem Israelem et transivit Iordanem venitque in Elam. Et direxerunt aciem Syri ex adverso David et pugnaverunt contra eum.
2SAM|10|18|Fugeruntque Syri a facie Israel; et occidit David de Syris septingentos currus et quadraginta milia peditum et Sobach principem militiae percussit, qui ibi mortuus est.
2SAM|10|19|Videntes autem universi reges, qui erant in praesidio Adadezer, se victos esse ab Israel, fecerunt pacem cum Israel et servierunt eis. Timueruntque Syri auxilium praebere ultra filiis Ammon.
2SAM|11|1|Factum est autem vertente anno, eo tempore quo solent reges ad bella procedere, misit David Ioab et servos suos cum eo et universum Israel, et vastaverunt filios Ammon et obsederunt Rabba; David autem remansit in Ierusalem.
2SAM|11|2|Et factum est vespere, ut surgeret David de strato suo et deambularet in solario domus regiae. Viditque de solario mulierem se lavantem; erat autem mulier pulchra valde.
2SAM|11|3|Misit ergo rex et requisivit quae esset mulier; nuntiatumque ei est quod ipsa esset Bethsabee filia Eliam uxor Uriae Hetthaei.
2SAM|11|4|Missis itaque David nuntiis, tulit eam; quae cum ingressa esset ad illum, dormivit cum ea, quae se sanctificaverat ab immunditia sua.
2SAM|11|5|Et reversa est domum suam; cum autem concepisset, mittens nuntiavit David et ait: " Concepi ".
2SAM|11|6|Misit autem David ad Ioab dicens: " Mitte ad me Uriam Hetthaeum ". Misitque Ioab Uriam ad David,
2SAM|11|7|et venit Urias ad David. Quaesivitque David quam recte ageret Ioab et populus, et quomodo administraretur bellum;
2SAM|11|8|et dixit David ad Uriam: " Descende in domum tuam et lava pedes tuos ". Et egressus est Urias de domo regis; secutusque est eum cibus regius.
2SAM|11|9|Dormivit autem Urias ante portam domus regiae cum aliis servis domini sui et non descendit ad domum suam.
2SAM|11|10|Nuntiatumque est David a dicentibus: " Non ivit Urias ad domum suam ". Et ait David ad Uriam: " Numquid non de via venisti? Quare non descendisti ad domum tuam? ".
2SAM|11|11|Et ait Urias ad David: " Arca et Israel et Iuda habitant in papilionibus, et dominus meus Ioab et servi domini mei super faciem terrae manent; et ego ingrediar domum meam, ut comedam et bibam et dormiam cum uxore mea? Per salutem tuam et per salutem animae tuae, non faciam rem hanc! ".
2SAM|11|12|Ait ergo David ad Uriam: " Mane hic etiam hodie, et cras dimittam te ". Mansit Urias in Ierusalem die illa et altera.
2SAM|11|13|Vocavit enim eum David, ut comederet coram se et biberet, et inebriavit eum. Qui egressus vespere dormivit in strato suo cum servis domini sui et in domum suam non descendit.
2SAM|11|14|Factum est ergo mane, et scripsit David epistulam ad Ioab misitque per manum Uriae
2SAM|11|15|scribens in epistula: " Ponite Uriam in prima acie, ubi fortissimum est proelium, et recedite ab eo, ut percussus intereat ".
2SAM|11|16|Igitur cum Ioab obsideret urbem, posuit Uriam in loco, quo sciebat viros esse fortissimos.
2SAM|11|17|Egressique viri de civitate bellabant adversum Ioab; et ceciderunt de populo, de servis David, et mortuus est etiam Urias Hetthaeus.
2SAM|11|18|Misit itaque Ioab et nuntiavit David omnia de proelio;
2SAM|11|19|praecepitque nuntio dicens: " Cum compleveris universos sermones proelii ad regem,
2SAM|11|20|si eum videris indignari et dixerit: "Quare accessistis ad urbem, ut proeliaremini? An ignorabatis quod desuper ex muro tela mittantur?
2SAM|11|21|Quis percussit Abimelech filium Ierobbaal? Nonne mulier misit super eum molam versatilem de muro, et mortuus est in Thebes? Quare iuxta murum accessistis?", dices: Etiam servus tuus Urias Hetthaeus occubuit ".
2SAM|11|22|Abiit ergo nuntius et venit et narravit David omnia, quae ei praeceperat Ioab.
2SAM|11|23|Et dixit nuntius ad David: " Quia praevaluerunt adversum nos viri et egressi sunt ad nos in agrum, nos, facto impetu, persecuti eos sumus usque ad portam civitatis.
2SAM|11|24|Et direxerunt iacula sagittarii ad servos tuos ex muro desuper; mortuique sunt de servis regis, quin etiam servus tuus Urias Hetthaeus mortuus est ".
2SAM|11|25|Et dixit David ad nuntium: " Haec dices Ioab: Non te affligat ista res; varius enim eventus est belli, et nunc hunc, nunc illum consumit gladius; corrobora proelium tuum adversus urbem, ut destruas eam. Et tu conforta eum ".
2SAM|11|26|Audivit autem uxor Uriae quod mortuus esset Urias vir suus et planxit eum.
2SAM|11|27|Transactoque luctu, misit David et introduxit eam domum suam, et facta est ei uxor peperitque ei filium. Et displicuit, quod fecerat David, coram Domino.
2SAM|12|1|Misit ergo Dominus Nathan ad David. Qui cum venisset ad eum, dixit ei: " Duo viri erant in civitate una, unus dives et alter pauper.
2SAM|12|2|Dives habebat oves et boves plurimos valde.
2SAM|12|3|Pauper autem nihil habebat omnino praeter ovem unam parvulam, quam emerat et nutrierat, et quae creverat apud eum cum filiis eius simul de pane illius comedens et de calice eius bibens et in sinu illius dormiens; eratque illi sicut filia.
2SAM|12|4|Cum autem peregrinus quidam venisset ad divitem, parcens ille sumere de ovibus et de bobus suis, ut exhiberet convivium peregrino illi, qui venerat ad se, tulit ovem viri pauperis et praeparavit cibos homini, qui venerat ad se ".
2SAM|12|5|Iratus autem indignatione David adversus hominem illum nimis dixit ad Nathan: " Vivit Dominus, quoniam filius mortis est vir, qui fecit hoc;
2SAM|12|6|ovem reddet in quadruplum, eo quod fecerit istud et non pepercerit ".
2SAM|12|7|Dixit autem Nathan ad David: " Tu es ille vir! Haec dicit Dominus, Deus Israel: Ego unxi te in regem super Israel et ego erui te de manu Saul;
2SAM|12|8|et dedi tibi domum domini tui et uxores domini tui in sinu tuo dedique tibi domum Israel et Iudae et, si parva sunt ista, adiciam tibi multo maiora.
2SAM|12|9|Quare ergo contempsisti verbum Domini, ut faceres malum in conspectu eius? Uriam Hetthaeum percussisti gladio et uxorem illius accepisti uxorem tibi et interfecisti eum gladio filiorum Ammon.
2SAM|12|10|Quam ob rem non recedet gladius de domo tua usque in sempiternum, eo quod despexeris me et tuleris uxorem Uriae Hetthaei, ut esset uxor tua.
2SAM|12|11|Itaque haec dicit Dominus: Ecce ego suscitabo super te malum de domo tua et tollam uxores tuas in oculis tuis et dabo proximo tuo, et dormiet cum uxoribus tuis in oculis solis huius.
2SAM|12|12|Tu enim fecisti abscondite; ego vero faciam istud in conspectu omnis Israel et in conspectu solis ".
2SAM|12|13|Et dixit David ad Nathan: " Peccavi Domino ". Dixitque Nathan ad David: Dominus quoque transtulit peccatum tuum; non morieris.
2SAM|12|14|Verumtamen quoniam blasphemare fecisti inimicos Domini propter hoc, filius, qui natus est tibi, morte morietur ".
2SAM|12|15|Et reversus est Nathan domum suam.Percussitque Dominus parvulum, quem peperat uxor Uriae David, et graviter aegrotavit;
2SAM|12|16|deprecatusque est David Dominum pro parvulo et ieiunavit David ieiunio et ingressus domum pernoctabat iacens super terram.
2SAM|12|17|Steterunt autem seniores domus eius iuxta eum cogentes eum, ut surgeret de terra; qui noluit neque comedit cum eis cibum.
2SAM|12|18|Accidit autem die septima, ut moreretur infans. Timueruntque servi David nuntiare ei quod mortuus esset parvulus; dixerunt enim: " Ecce, cum parvulus adhuc viveret, loquebamur ad eum, et non audiebat vocem nostram. Nunc quomodo dicemus: "Mortuus est puer"? Peius patrabit! ".
2SAM|12|19|Cum ergo vidisset David servos suos mussitantes, intellexit quod mortuus esset infantulus dixitque ad servos suos: " Num mortuus est puer?. Qui responderunt ei: " Mortuus est ".
2SAM|12|20|Surrexit igitur David de terra et lotus unctusque est; cumque mutasset vestem, ingressus est domum Domini et adoravit et venit in domum suam petivitque, ut ponerent ei panem, et comedit.
2SAM|12|21|Dixerunt autem ei servi sui: " Quid est quod fecisti? Propter infantem, cum adhuc viveret, ieiunasti et flebas; mortuo autem puero, surrexisti et comedisti panem ".
2SAM|12|22|Qui ait: " Propter infantem, dum adhuc viveret, ieiunavi et flevi. Dicebam enim: Quis scit, si forte miserebitur mei Dominus, et vivet infans?
2SAM|12|23|Nunc autem, quia mortuus est, quare ieiuno? Numquid potero revocare eum amplius? Ego vadam magis ad eum, ille vero non revertetur ad me ".
2SAM|12|24|Et consolatus est David Bethsabee uxorem suam ingressusque ad eam dormivit cum ea, quae genuit filium; et vocavit nomen eius Salomon. Et Dominus dilexit eum
2SAM|12|25|misitque in manu Nathan prophetae et vocavit nomen eius Iedidia (id est Amabilis Domino) propter Dominum.
2SAM|12|26|Igitur pugnavit Ioab contra Rabba filiorum Ammon et expugnavit urbem regiam.
2SAM|12|27|Misitque Ioab nuntios ad David dicens: " Dimicavi adversum Rabba et cepi urbem aquarum;
2SAM|12|28|nunc igitur congrega reliquam partem populi et obside civitatem et cape eam, ne, cum a me capta fuerit urbs, nomine meo vocetur ".
2SAM|12|29|Congregavit itaque David omnem populum et profectus est adversum Rabba; cumque dimicasset, cepit eam.
2SAM|12|30|Et tulit diadema Melchom de capite eius, pondo auri talentum, habens gemmam pretiosissimam, quod venit super caput David. Sed et praedam civitatis asportavit multam valde,
2SAM|12|31|populum quoque eius educens condemnavit ad operam lapicidinarum et ad secures et dolabras ferreas et transtulit eos ad opus laterum; sic fecit universis civitatibus filiorum Ammon. Et reversus est David et omnis exercitus Ierusalem.
2SAM|13|1|Factum est autem post haec, ut Absalom filii David soro rem speciosissimam, vocabulo Thamar, adamaret Amnon filius David.
2SAM|13|2|Et angustiatus est Amnon, ita ut aegrotaret propter amorem Thamar sororis suae, quia, cum esset virgo, difficile ei videbatur ut quippiam inhoneste ageret cum ea.
2SAM|13|3|Erat autem Amnonis amicus nomine Ionadab filius Samma fratris David, vir callidus valde.
2SAM|13|4|Qui dixit ad eum: " Quare sic attenuaris macie, fili regis, per singulos dies? Cur non indicas mihi? ". Dixitque ei Amnon: " Thamar sororem Absalom fratris mei amo ".
2SAM|13|5|Cui respondit Ionadab: " Cuba super lectulum tuum et languorem simula. Cumque venerit pater tuus, ut visitet te, dic ei: "Veniat, oro, Thamar soror mea, ut det mihi cibum et faciat in oculis meis pulmentum, ut videam et comedam de manu eius" ".
2SAM|13|6|Accubuit itaque Amnon et simulavit languorem. Cumque venisset rex ad visitandum eum, ait Amnon ad regem: " Veniat, obsecro, Thamar soror mea, ut faciat in oculis meis duas sorbitiunculas, et cibum capiam de manu eius.
2SAM|13|7|Misit ergo David ad Thamar domum dicens: " Veni in domum Amnon fratris tui et fac ei pulmentum ".
2SAM|13|8|Venitque Thamar in domum Amnon fratris sui; ille autem iacebat. Quae tollens farinam commiscuit et conficiens in oculis eius coxit sorbitiunculas.
2SAM|13|9|Tollensque sartaginem effudit, quod coxerat, et posuit coram eo. Noluit comedere; dixitque Amnon: " Eicite universos a me ". Cumque exissent omnes,
2SAM|13|10|dixit Amnon ad Thamar: " Infer cibum in conclave, ut vescar de manu tua. Tulit ergo Thamar sorbitiunculas, quas fecerat, et intulit ad Amnon fratrem suum in conclave.
2SAM|13|11|Cumque obtulisset ei cibum, apprehendit eam et ait: " Veni, cuba mecum, soror mea ".
2SAM|13|12|Quae respondit ei: " Noli, frater mi, noli opprimere me! Neque enim hoc fas est in Israel; noli facere stultitiam hanc.
2SAM|13|13|Et ego quo ibo in opprobrio meo? Et tu eris quasi unus de insipientibus in Israel; quin potius loquere ad regem, et non negabit me tibi ".
2SAM|13|14|Noluit autem acquiescere precibus eius, sed praevalens viribus oppressit eam et cubavit cum illa.
2SAM|13|15|Et exosam eam habuit Amnon magno odio nimis, ita ut maius esset odium, quo oderat eam, amore, quo ante dilexerat. Dixitque ei Amnon: " Surge, vade! ".
2SAM|13|16|Quae respondit ei: " Ne fiat, frater mi, quia maius est hoc malum, quod nunc agis adversum me expellens me, quam quod ante fecisti ". Et noluit audire eam;
2SAM|13|17|sed vocato puero, qui ministrabat ei, dixit: " Eice hanc a me foras et claude ostium post eam ".
2SAM|13|18|Quae induta erat talari tunica; huiusmodi enim filiae regis virgines palliis vestibus utebantur. Eiecit itaque eam minister illius foras clausitque fores post eam.
2SAM|13|19|Quae aspergens pulverem capiti suo, scissa talari tunica impositisque manibus super caput suum, ibat ingrediens et clamans.
2SAM|13|20|Dixit autem ei Absalom frater suus: " Num Amnon frater tuus fuit tecum? Sed nunc, soror, tace: frater tuus est; neque affligas cor tuum pro re hac. Mansit itaque Thamar desolata in domo Absalom fratris sui.
2SAM|13|21|Cum autem audisset rex David omnia haec, iratus est valde; et noluit contristare spiritum Amnon filii sui, quoniam diligebat eum, quia primogenitus erat ei.
2SAM|13|22|Porro non est locutus Absalom ad Amnon nec malum nec bonum; oderat enim Absalom Amnon, eo quod violasset Thamar sororem suam.
2SAM|13|23|Factum est autem post tempus biennii, ut tonderentur oves Absalom in Baalhasor, quae est iuxta Ephraim; et vocavit Absalom omnes filios regis.
2SAM|13|24|Venitque ad regem et ait ad eum: " Ecce tondentur oves servi tui; veniat, oro, rex cum servis suis ad servum tuum ".
2SAM|13|25|Dixitque rex ad Absalom: " Noli, fili mi, noli rogare, ut veniamus omnes et gravemus te ". Cum autem cogeret eum, et noluisset ire, benedixit ei.
2SAM|13|26|Et ait Absalom: " Si non vis venire, veniat, obsecro, nobiscum saltem Amnon frater meus ". Dixitque ad eum rex: " Cur vadet tecum? ".
2SAM|13|27|Coegit itaque eum Absalom, et dimisit cum eo Amnon et universos filios regis.Fecitque Absalom convivium quasi convivium regis.
2SAM|13|28|Praecepit autem Absalom pueris suis dicens: " Observate. Cum hilarior fuerit Amnon vino, et dixero vobis: Percutite Amnon et interficite eum!, nolite timere; ego enim sum, qui praecepi vobis. Roboramini et estote viri fortes ".
2SAM|13|29|Fecerunt ergo pueri Absalom adversum Amnon, sicut praeceperat eis Absalom; surgentesque omnes filii regis ascenderunt singuli mulos suos et fugerunt.
2SAM|13|30|Cumque adhuc pergerent in itinere, fama praevenit ad David dicens: " Percussit Absalom omnes filios regis, et non remansit ex eis saltem unus.
2SAM|13|31|Surrexit itaque rex et scidit vestimenta sua et prostravit se super terram; et omnes servi ipsius, qui assistebant ei, sciderunt vestimenta sua.
2SAM|13|32|Respondens autem Ionadab filius Samma fratris David dixit: " Ne aestimet dominus meus quod omnes pueri filii regis occisi sint; Amnon solus mortuus est, quoniam in ore Absalom hoc erat positum ex die, qua oppressit Thamar sororem eius.
2SAM|13|33|Nunc ergo ne ponat dominus meus rex super cor suum verbum istud dicens: Omnes filii regis occisi sunt", quoniam Amnon solus mortuus est ".
2SAM|13|34|Fugit autem Absalom.Et levavit puer speculator oculos suos et aspexit, et ecce populus multus veniebat per viam Oronaim ex latere montis in descensu; et venit speculator et nuntiavit regi dicens: " Video homines per viam Oronaim ".
2SAM|13|35|Dixit autem Ionadab ad regem: " Ecce filii regis adsunt! Iuxta verbum servi tui sic factum est ".
2SAM|13|36|Cumque cessasset loqui, apparuerunt et filii regis et intrantes levaverunt vocem suam et fleverunt; sed et rex et omnes servi eius fleverunt ploratu magno nimis.
2SAM|13|37|Porro Absalom fugiens abiit ad Tholmai filium Ammiud regem Gesur. Luxit ergo David filium suum cunctis diebus.
2SAM|13|38|Absalom autem, cum fugisset et venisset in Gesur, fuit ibi tribus annis.
2SAM|13|39|Cessavitque spiritus regis adversari Absalom, eo quod consolatus esset super Amnon interitu.
2SAM|14|1|Intellegens autem Ioab filius Sarviae quod cor regis ver sum esset ad Absalom,
2SAM|14|2|misit Thecuam et tulit inde mulierem sapientem dixitque ad eam: " Lugere te simula et induere veste lugubri et ne ungaris oleo, ut sis quasi mulier plurimo iam tempore lugens mortuum.
2SAM|14|3|Et ingredieris ad regem et loqueris ad eum sermones huiuscemodi ". Posuit autem Ioab verba in ore eius.
2SAM|14|4|Itaque, cum ingressa fuisset mulier Thecuites ad regem, cecidit coram eo super terram et adoravit et dixit: " Serva me, rex ".
2SAM|14|5|Et ait ad eam rex: " Quid causae habes? ". Quae respondit: " Heu, mulier vidua ego sum: mortuus est vir meus.
2SAM|14|6|Et ancillae tuae erant duo filii, qui rixati sunt adversum se in agro, nullusque erat, qui eos interveniens prohibere posset; et percussit alter alterum et interfecit eum.
2SAM|14|7|Et ecce consurgens universa cognatio adversum ancillam tuam dicit: Trade eum, qui percussit fratrem suum, ut occidamus eum pro anima fratris sui, quem interfecit, et deleamus heredem". Et quaerunt exstinguere scintillam meam, quae relicta est, ut non supersit viro meo nomen et reliquiae super terram ".
2SAM|14|8|Et ait rex ad mulierem: " Vade in domum tuam, et ego iubebo de te ".
2SAM|14|9|Dixitque mulier Thecuites ad regem: " In me, domine mi rex, iniquitas et in domum patris mei; rex autem et thronus eius sit innocens ".
2SAM|14|10|Et ait rex: " Qui contradixerit tibi, adduc eum ad me, et ultra non addet ut tangat te ".
2SAM|14|11|Quae ait: " Recordetur rex Domini Dei sui, ut non augeat ultor sanguinis perniciem, et nequaquam interficiant filium meum ". Qui ait: " Vivit Dominus, quia non cadet de capillis filii tui super terram ".
2SAM|14|12|Dixit ergo mulier: " Loquatur ancilla tua ad dominum meum regem verbum. Et ait: " Loquere ".
2SAM|14|13|Dixitque mulier: " Quare cogitasti istiusmodi rem contra populum Dei? Eo enim quod rex locutus est verbum istud, hoc est quasi delictum, quia rex noluit reducere eiectum suum.
2SAM|14|14|Omnes morimur et quasi aquae sumus, quae delabuntur in terram, quae non colliguntur; nec tamen vult perire Deus animam, sed retractat cogitans, ne penitus pereat, qui abiectus est.
2SAM|14|15|Nunc igitur veni, ut loquar ad regem dominum meum verbum hoc, quia populus terruit me. Et dixit ancilla tua: Loquar ad regem, si quo modo faciat rex verbum ancillae suae.
2SAM|14|16|Nam audiet rex, ut liberet ancillam suam de manu illius, qui vult delere me et filium meum simul de hereditate Dei.
2SAM|14|17|Dixit ergo ancilla tua: Fiat verbum domini mei regis mihi in quietem. Sicut enim angelus Dei, sic est dominus meus rex, ut audiat et discernat bonum et malum. Et Dominus Deus tuus sit tecum! ".
2SAM|14|18|Et respondens rex dixit ad mulierem: " Ne abscondas a me verbum, quod te interrogo ". Dixitque mulier: " Loquatur dominus meus rex ".
2SAM|14|19|Et ait rex: " Numquid manus Ioab tecum est in omnibus istis? ". Respondit mulier et ait: " Per salutem animae tuae, domine mi rex, nec ad dextram nec ad sinistram potest deviari ab omnibus his, quae locutus est dominus meus rex; servus enim tuus Ioab ipse praecepit mihi et ipse posuit in os ancillae tuae omnia verba haec;
2SAM|14|20|ut verterem figuram rei huius, servus tuus Ioab fecit istud. Tu autem, domine mi, sapiens es, sicut habet sapientiam angelus Dei, ut intellegas omnia, quae fiunt super terram ".
2SAM|14|21|Et ait rex ad Ioab: " Ecce hoc facio; vade igitur et revoca puerum Absalom ".
2SAM|14|22|Cadensque Ioab super faciem suam in terram adoravit et benedixit regi. Et dixit Ioab: " Hodie intellexit servus tuus quia inveni gratiam in oculis tuis, domine mi rex; fecisti enim sermonem servi tui ".
2SAM|14|23|Surrexit ergo Ioab et abiit in Gesur et adduxit Absalom in Ierusalem.
2SAM|14|24|Dixit autem rex: " Revertatur in domum suam et faciem meam non videat. Reversus est itaque Absalom in domum suam et faciem regis non vidit.
2SAM|14|25|Porro sicut Absalom vir non erat pulcher in omni Israel, qui valde laudaretur, a vestigio pedis usque ad verticem non erat in eo ulla macula.
2SAM|14|26|Et quando tondebatur capillus - semel autem in anno tondebatur, quia gravabat eum caesaries - ponderabat capillos capitis sui ducentis siclis pondere regio.
2SAM|14|27|Nati sunt autem Absalom filii tres et filia una, nomine Thamar, eleganti forma.
2SAM|14|28|Mansitque Absalom Ierusalem duobus annis et faciem regis non vidit.
2SAM|14|29|Misit itaque ad Ioab, ut mitteret eum ad regem; qui noluit venire ad eum. Cumque secundo misisset, et ille noluisset venire,
2SAM|14|30|dixit servis suis: " Videte agrum Ioab iuxta agrum meum habentem messem hordei; ite igitur et succendite eum igni ". Succenderunt ergo servi Absalom segetem igni. Et venientes servi Ioab, scissis vestibus suis, dixerunt: " Succenderunt servi Absalom agrum igni! ".
2SAM|14|31|Surrexitque Ioab et venit ad Absalom in domum eius et dixit: " Quare succenderunt servi tui segetem meam igni? ".
2SAM|14|32|Et respondit Absalom ad Ioab: " Misi ad te obsecrans, ut venires ad me, et mitterem te ad regem, ut diceres ei: "Quare veni de Gesur? Melius mihi erat adhuc ibi esse". Obsecro ergo, ut videam faciem regis; quod si est in me iniquitas, interficiat me ".
2SAM|14|33|Ingressus Ioab ad regem nuntiavit ei. Vocatusque Absalom intravit ad regem et adoravit super faciem in terra coram eo; osculatusque est rex Absalom.
2SAM|15|1|Post haec fecit sibi Absalom currus et equos et quinqua ginta viros, qui praecederent eum.
2SAM|15|2|Et mane consurgens Absalom stabat iuxta viam portae; et omnem virum, qui habebat negotium, ut veniret ad regis iudicium, vocabat Absalom ad se et dicebat: " De qua civitate es tu? ". Qui respondens aiebat: " Ex una tribu Israel ego sum servus tuus ".
2SAM|15|3|Respondebatque ei Absalom: " Vide, sermones tui sunt boni et iusti, sed non est qui te audiat constitutus a rege ". Dicebatque Absalom:
2SAM|15|4|" Quis me constituat iudicem in terra, ut ad me veniant omnes, qui habent negotium iudicandum, et iustificem eos? ".
2SAM|15|5|Sed et cum accederet ad eum homo, ut se prostraret coram illo, extendebat manum suam et apprehendens osculabatur eum.
2SAM|15|6|Faciebatque hoc omni Israel, qui veniebat ad iudicium, ut audiretur a rege, et sollicitabat corda virorum Israel.
2SAM|15|7|Post quattuor autem annos dixit Absalom ad regem: " Vadam, quaeso, et reddam in Hebron vota mea, quae vovi Domino.
2SAM|15|8|Votum enim vovit servus tuus, cum esset in Gesur Syriae, dicens: Si reduxerit me Dominus in Ierusalem, sacrificabo Domino ".
2SAM|15|9|Dixitque ei rex. " Vade in pace ". Et surrexit et abiit in Hebron.
2SAM|15|10|Misit autem Absalom exploratores in universas tribus Israel dicens: " Statim ut audieritis clangorem bucinae, dicite: "Factus est rex Absalom in Hebron" ".
2SAM|15|11|Porro cum Absalom ierunt ducenti viri de Ierusalem vocati, euntes simplici corde et causam penitus ignorantes.
2SAM|15|12|Accersivit quoque Absalom, cum immolaret victimas, Achitophel Gilonitem consiliarium David de civitate sua Gilo. Et facta est coniuratio valida; populusque concurrens augebatur cum Absalom.
2SAM|15|13|Venit igitur nuntius ad David dicens: " Toto corde universus Israel sequitur Absalom ".
2SAM|15|14|Et ait David servis suis, qui erant cum eo in Ierusalem: " Surgite, fugiamus; neque enim erit nobis effugium a facie Absalom. Festinate egredi, ne festinans occupet nos et impellat super nos ruinam et percutiat civitatem in ore gladii ".
2SAM|15|15|Dixeruntque servi regis ad eum: " In omnibus, quaecumque elegerit dominus noster rex, ecce servi tui sumus ".
2SAM|15|16|Egressus est ergo rex et universa domus eius post eum et dereliquit rex decem mulieres concubinas ad custodiendam domum.
2SAM|15|17|Egressusque rex et omnis populus post eum steterunt ad ultimam domum.
2SAM|15|18|Et universi servi eius transierunt iuxta eum; et omnes Cherethi et Phelethi et omnes Getthaei, sescenti viri, qui secuti eum fuerant de Geth, transierunt coram rege.
2SAM|15|19|Dixit autem rex ad Ethai Getthaeum: " Cur venis etiam tu nobiscum? Revertere et habita cum rege, quia alienigena es, immo et exsul de loco tuo.
2SAM|15|20|Heri venisti, et hodie compellam te vagari nobiscum, cum ego vadam, quo iturus sum? Revertere et reduc tecum fratres tuos, et Dominus faciat tecum misericordiam et veritatem ".
2SAM|15|21|Et respondit Ethai regi dicens: " Vivit Dominus et vivit dominus meus rex, in quocumque loco fuerit dominus meus rex, sive ad mortem sive ad vitam, ibi erit servus tuus ".
2SAM|15|22|Et ait David Ethai: " Veni et transi ". Et transivit Ethai Getthaeus et omnes viri eius et omnes parvuli, qui cum eo erant.
2SAM|15|23|Omnisque terra flebat voce magna, et universus populus transibat. Rex quoque transgrediebatur torrentem Cedron, et cunctus populus incedebat contra viam deserti.
2SAM|15|24|Venit autem et Sadoc et universi Levitae cum eo portantes arcam foederis Dei; et deposuerunt arcam Dei. Et sacrificavit Abiathar, donec omnis populus egressus fuerat de civitate.
2SAM|15|25|Et dixit rex ad Sadoc: " Reporta arcam Dei in urbem. Si invenero gratiam in oculis Domini, reducet me et ostendet mihi eam et habitationem suam.
2SAM|15|26|Si autem dixerit: "Non places mihi", praesto sum: faciat, quod bonum est coram se ".
2SAM|15|27|Et dixit rex ad Sadoc sacerdotem: " Videsne? Revertere in civitatem in pace; et Achimaas filius tuus et Ionathan filius Abiathar, duo filii vestri sint vobiscum.
2SAM|15|28|Ecce ego morabor ad vada deserti, donec veniat sermo a vobis indicans mihi ".
2SAM|15|29|Reportaverunt igitur Sadoc et Abiathar arcam Dei Ierusalem et manserunt ibi.
2SAM|15|30|Porro David ascendebat clivum Olivarum scandens et flens, operto capite et nudis pedibus incedens; sed et omnis populus, qui erat cum eo, operto capite ascendebat plorans.
2SAM|15|31|Nuntiatum est autem David quod et Achitophel esset in coniuratione cum Absalom; dixitque David: " Infatua, quaeso, Domine, consilium Achitophel.
2SAM|15|32|Cumque ascendisset David summitatem montis, in quo adorabatur Deus, ecce occurrit ei Chusai Arachites, scissa veste et terra pleno capite.
2SAM|15|33|Et dixit ei David: " Si veneris mecum, eris mihi oneri;
2SAM|15|34|Si autem in civitatem revertaris et dixeris Absalom: "Servus tuus ego, rex, ero; servus patris tui ego fui prius, nunc autem ego sum servus tuus", dissipabis mihi consilium Achitophel.
2SAM|15|35|Habes autem tecum Sadoc et Abiathar sacerdotes; et omne verbum, quodcumque audieris de domo regis, indicabis Sadoc et Abiathar sacerdotibus.
2SAM|15|36|Sunt autem cum eis duo filii eorum: Achimaas Sadoc et Ionathan Abiathar; et mittetis per eos ad me omne verbum, quod audieritis ".
2SAM|15|37|Veniente ergo Chusai amico David in civitatem, Absalom quoque ingressus est Ierusalem.
2SAM|16|1|Cumque David transisset paululum montis verticem, apparuit Siba puer Meribbaal in occursum eius cum duobus asinis stratis, qui onerati erant ducentis panibus et centum alligaturis uvae passae et centum fasciculis fructuum aestivorum et utre vini.
2SAM|16|2|Et dixit rex Sibae: " Quid sibi volunt haec? ". Responditque Siba: " Asini domesticis regis ad sedendum; et panes et fructus aestivi ad vescendum pueris tuis; vinum autem, ut bibat, si quis defecerit in deserto.
2SAM|16|3|Et ait rex: " Ubi est filius domini tui? ". Responditque Siba regi: " Remansit in Ierusalem dicens: "Hodie restituet mihi domus Israel regnum patris mei" ".
2SAM|16|4|Et ait rex Sibae: " Ecce, tua sint omnia, quae fuerunt Meribbaal ". Dixitque Siba: " Adoro; inveniam gratiam coram te, domine mi rex ".
2SAM|16|5|Venit ergo rex David usque Bahurim, et ecce egrediebatur inde vir de cognatione domus Saul nomine Semei filius Gera; procedebat egrediens et maledicens
2SAM|16|6|mittebatque lapides contra David et contra universos servos regis David. Omnis autem populus et universi viri fortissimi a dextro et sinistro latere regis incedebant.
2SAM|16|7|Ita autem loquebatur Semei, cum malediceret regi: " Egredere, egredere, vir sanguinum et vir Belial!
2SAM|16|8|Reddidit tibi Dominus universum sanguinem domus Saul, quoniam invasisti regnum eius; et dedit Dominus regnum in manu Absalom filii tui; et ecce premunt te mala tua, quoniam vir sanguinum es ".
2SAM|16|9|Dixit autem Abisai filius Sarviae regi: " Quare maledicit canis hic mortuus domino meo regi? Vadam et amputabo caput eius ".
2SAM|16|10|Et ait rex: "Quid mihi et vobis filii Sarviae? Si maledicit, et si Dominus praecepit ei, ut malediceret David, quis est qui audeat dicere: Quare sic fecisti?" ".
2SAM|16|11|Et ait rex Abisai et universis servis suis: " Ecce filius meus, qui egressus est de visceribus meis, quaerit animam meam; quanto magis nunc iste filius Beniaminita. Dimittite eum, ut maledicat iuxta praeceptum Domini.
2SAM|16|12|Fortasse respiciet Dominus afflictionem meam et reddet mihi bonum pro maledictione hac hodierna ".
2SAM|16|13|Ambulabat itaque David et socii eius per viam; Semei autem per iugum montis ex latere gradiebatur maledicens et mittens lapides adversum eum terramque spargens.
2SAM|16|14|Venit itaque rex et universus populus cum eo lassus usque ad aquas, et refocillati sunt ibi.
2SAM|16|15|Absalom autem et omnis populus eius, viri Israel, ingressi sunt Ierusalem, sed et Achitophel cum eo.
2SAM|16|16|Cum autem venisset Chusai Arachites amicus David ad Absalom, locutus est ad eum: " Vivat rex! Vivat rex! ".
2SAM|16|17|Ad quem Absalom: "Haec est, inquit, gratia tua ad amicum tuum? Quare non isti cum amico tuo? ".
2SAM|16|18|Responditque Chusai ad Absalom: " Nequaquam; quia, quem elegit Dominus, et hic populus et omnis Israel, illius ero et cum eo manebo.
2SAM|16|19|Sed, ut et hoc inferam, cui ego serviturus sum? Nonne filio regis? Sicut parui patri tuo, sic parebo et tibi ".
2SAM|16|20|Dixit autem Absalom ad Achitophel: " Inite consilium quid agere debeamus ".
2SAM|16|21|Et ait Achitophel ad Absalom: " Ingredere ad concubinas patris tui, quas dimisit ad custodiendam domum; ut, cum audierit omnis Israel quod foedaveris patrem tuum, roborentur manus omnium, qui tecum sunt ".
2SAM|16|22|Tetenderunt igitur Absalom tabernaculum in solario; ingressusque est ad concubinas patris sui coram universo Israel.
2SAM|16|23|Consilium autem Achitophel, quod dabat in diebus illis, quasi si quis consuleret Deum; sic erat omne consilium Achitophel, et cum esset cum David et cum esset cum Absalom.
2SAM|17|1|Dixitque Achitophel ad Ab salom: " Eligam mihi duode cim milia virorum et consurgens persequar David hac nocte
2SAM|17|2|et irruens super eum, quippe qui lassus est et solutis manibus, terrebo eum. Cumque fugerit omnis populus, qui cum eo est, percutiam regem desolatum
2SAM|17|3|et reducam universum populum ad te, sicut revertitur sponsa ad virum suum; unius solummodo viri animam quaeris, et omnis populus erit in pace.
2SAM|17|4|Placuitque sermo eius Absalom et cunctis maioribus natu Israel.
2SAM|17|5|Ait autem Absalom: " Vocate et Chusai Arachiten, et audiamus quid etiam ipse dicat ".
2SAM|17|6|Cumque venisset Chusai ad Absalom, ait Absalom ad eum: " Huiuscemodi sermonem locutus est Achitophel; verbum eius facere debemus an non? Tu loquere ".
2SAM|17|7|Et dixit Chusai ad Absalom: " Non bonum consilium, quod dedit Achitophel hac vice ".
2SAM|17|8|Et rursum intulit Chusai: " Tu nosti patrem tuum et viros, qui cum eo sunt, esse fortissimos et amaro animo, veluti ursa in saltu catulis orbata; sed et pater tuus vir bellator est nec morabitur cum populo:
2SAM|17|9|ecce nunc latitat in aliqua fovea aut in aliquo alio loco. Et, cum ceciderit unus quilibet in principio, certo audient et dicent: "Facta est plaga in populo, qui sequitur Absalom".
2SAM|17|10|Et fortissimus quoque, cuius cor est quasi leonis, pavore solvetur; scit enim omnis Israel fortem esse patrem tuum et robustos omnes, qui cum eo sunt.
2SAM|17|11|Sed hoc mihi videtur rectum esse consilium: congregetur ad te universus Israel a Dan usque Bersabee, quasi arena maris innumerabilis, et tu ipse gradieris in proelium;
2SAM|17|12|et irruemus super eum, in quocumque loco fuerit inventus, et operiemus eum sicut cadere solet ros super terram; et non remanebit de eo et de omnibus viris, qui cum eo sunt, ne unus quidem.
2SAM|17|13|Quod si urbem aliquam fuerit ingressus, applicabit omnis Israel civitati illi funes, et trahemus eam in torrentem, ut non reperiatur nec calculus quidem ex ea ".
2SAM|17|14|Dixitque Absalom et omnis vir Israel: " Melius consilium Chusai Arachitae consilio Achitophel ". Dominus enim statuerat dissipare consilium Achitophel utile, ut induceret Dominus super Absalom malum.
2SAM|17|15|Et ait Chusai Sadoc et Abiathar sacerdotibus: " Hoc et hoc modo consilium dedit Achitophel Absalom et senibus Israel, et ego tale et tale dedi consilium;
2SAM|17|16|nunc ergo mittite cito et nuntiate David dicentes: "Ne moreris nocte hac ad vada deserti, sed absque dilatione transgredere, ne absorbeatur rex et omnis populus, qui cum eo est" ".
2SAM|17|17|Ionathan autem et Achimaas stabant iuxta fontem Rogel; abiit ancilla et nuntiavit eis, et illi profecti sunt, ut referrent ad regem David nuntium; non enim poterant introire civitatem, ne viderentur.
2SAM|17|18|Vidit autem eos quidam iuvenis et indicavit Absalom; illi vero concito gradu profecti ingressi sunt domum cuiusdam viri in Bahurim, qui habebat puteum in vestibulo suo, et descenderunt in eum.
2SAM|17|19|Tulit autem mulier et expandit velamen super os putei et sparsit super illud ptisanas, et sic res latuit.
2SAM|17|20|Cumque venissent servi Absalom ad mulierem in domum, dixerunt: " Ubi est Achimaas et Ionathan? ". Et respondit eis mulier: " Transierunt hinc ad aquas ". At hi, qui quaerebant, cum non repperissent, reversi sunt Ierusalem.
2SAM|17|21|Cumque abissent, ascenderunt illi de puteo et pergentes nuntiaverunt regi David atque dixerunt: " Surgite et transite cito fluvium, quoniam huiuscemodi dedit consilium contra vos Achitophel ".
2SAM|17|22|Surrexit ergo David et omnis populus, qui erat cum eo, et transierunt Iordanem, donec dilucesceret; et ne unus quidem residuus fuit, qui non transisset fluvium.
2SAM|17|23|Porro Achitophel videns quod non fuisset factum consilium suum, stravit asinum suum et surrexit et abiit in domum suam in civitatem suam et, disposita domo sua, laqueo se suspendit et interiit; et sepultus est in sepulcro patris sui.
2SAM|17|24|David autem venit in Mahanaim, et Absalom transivit Iordanem, ipse et omnis vir Israel cum eo.
2SAM|17|25|Amasam vero constituerat Absalom pro Ioab super exercitum; Amasa autem erat filius viri, qui vocabatur Iether Ismaelites, qui ingressus est ad Abigail filiam Isai sororem Sarviae, quae fuit mater Ioab.
2SAM|17|26|Et castrametatus est Israel cum Absalom in terra Galaad.
2SAM|17|27|Cumque venisset David in Mahanaim, Sobi filius Naas de Rabba filiorum Ammon et Machir filius Ammiel de Lodabar et Berzellai Galaadites de Rogelim
2SAM|17|28|obtulerunt ei stratoria et tapetia et pelves et vasa fictilia, frumentum et hordeum et farinam, frixum cicer et fabam et lentem
2SAM|17|29|et mel et butyrum, oves et pingues vitulos; dederuntque David et populo, qui cum eo erat, ad vescendum; suspicati enim sunt populum fame et siti fuisse fatigatum in deserto.
2SAM|18|1|Igitur, recensito David populo suo, constituit super eum tribunos et centuriones.
2SAM|18|2|Et divisit David populum in tres partes: tertiam partem sub manu Ioab et tertiam sub manu Abisai filii Sarviae fratris Ioab et tertiam in manu Ethai, qui erat de Geth. Dixitque rex ad populum: " Egrediar et ego vobiscum ".
2SAM|18|3|Et respondit populus: " Non exibis. Sive enim fugerimus, non magnopere ad eos de nobis pertinebit; et si media pars ceciderit e nobis, non satis curabunt, sed tu unus pro decem milibus computaris. Melius est igitur, ut sis nobis ex urbe praesidio ".
2SAM|18|4|Ad quos rex ait: " Quod vobis rectum videtur, hoc faciam ". Stetit ergo rex iuxta portam; egrediebaturque populus per turmas suas centeni et milleni.
2SAM|18|5|Et praecepit rex Ioab et Abisai et Ethai dicens: " Leniter mihi agite cum puero Absalom ". Et omnis populus audiebat praecipientem regem cunctis principibus pro Absalom.
2SAM|18|6|Itaque egressus est populus in campum contra Israel, et factum est proelium in saltu Ephraim.
2SAM|18|7|Et caesus est ibi populus Israel ab exercitu David; factaque est ibi plaga magna in die illa viginti milium hominum.
2SAM|18|8|Fuit autem ibi proelium dispersum super faciem omnis terrae; et multo plures erant, quos saltus consumpserat de populo, quam hi, quos voraverat gladius in die illa.
2SAM|18|9|Accidit autem, ut occurreret Absalom servis David sedens mulo; cumque ingressus fuisset mulus subter condensam quercum et magnam, adhaesit caput eius quercui, et mansit suspensus inter caelum et terram; mulus, cui insederat, pertransivit.
2SAM|18|10|Vidit autem hoc quispiam et nuntiavit Ioab dicens: " Vidi Absalom pendere de quercu ".
2SAM|18|11|Et ait Ioab viro, qui nuntiaverat ei: " Si vidisti, quare non confodisti eum in terra? Ego vero dedissem tibi decem argenti siclos et unum balteum ".
2SAM|18|12|Qui dixit ad Ioab: " Et si appenderes in manibus meis mille argenteos, nequaquam mitterem manum meam in filium regis. Audientibus enim nobis, praecepit rex tibi et Abisai et Ethai dicens: "Custodite, quisquis sit, puerum Absalom!".
2SAM|18|13|Sed et si fecissem contra animam meam infideliter, nequaquam hoc regem latere potuisset, et tu stares ex adverso ".
2SAM|18|14|Et ait Ioab: " Non ita praestolabor coram te ". Tulit ergo tres lanceas in manu sua et infixit eas in corde Absalom, cum adhuc palpitaret haerens in quercu;
2SAM|18|15|et cucurrerunt decem iuvenes armigeri Ioab et percutientes interfecerunt eum.
2SAM|18|16|Cecinit autem Ioab bucina, et destitit populus persequi fugientem Israel, quia Ioab retinuit populum.
2SAM|18|17|Et tulerunt Absalom et proiecerunt eum in saltu in foveam grandem et erexerunt super eum acervum lapidum magnum nimis; omnis autem Israel fugit in tabernacula sua.
2SAM|18|18|Porro Absalom erexerat sibi, cum adhuc viveret, lapidem, qui est in valle Regis; dixerat enim: " Non habeo filium, qui memoriam servabit nominis mei ". Vocavitque titulum nomine suo, et appellatur Manus Absalom usque ad hanc diem.
2SAM|18|19|Achimaas autem filius Sadoc ait: " Curram et nuntiabo regi, quia iudicium fecerit ei Dominus de manu inimicorum eius ".
2SAM|18|20|Ad quem Ioab dixit: " Non es vir boni nuntii in hac die, sed nuntiabis in alia; hodie enim non nuntiabis bona, eo quod filius regis est mortuus.
2SAM|18|21|Et ait Ioab Aethiopi: " Vade et nuntia regi, quae vidisti ". Adoravit Aethiops Ioab et cucurrit.
2SAM|18|22|Rursus autem Achimaas filius Sadoc dixit ad Ioab: " Quidquid evenerit, etiam ego curram post Aethiopem! ". Dixitque Ioab: " Quid vis currere, fili mi? Non erit tibi merces pro bono nuntio ".
2SAM|18|23|Qui respondit: " Quidquid evenerit, curram ". Et ait ei: " Curre! ". Currens ergo Achimaas per viam regionis transivit Aethiopem.
2SAM|18|24|David autem sedebat inter duas portas; speculator vero, qui ierat in solarium portae super murum, elevans oculos vidit hominem currentem solum
2SAM|18|25|et exclamans indicavit regi. Dixitque rex: " Si solus est, bonus est nuntius in ore eius ". Properante autem illo et accedente propius,
2SAM|18|26|vidit speculator hominem alterum currentem, et clamavit speculator ad ianitorem: " Apparet mihi homo currens solus ". Dixitque rex: " Et iste bonus est nuntius ".
2SAM|18|27|Speculator autem: " Contemplor, ait, cursum prioris quasi cursum Achimaas filii Sadoc ". Et ait rex: " Vir bonus est et nuntium portans bonum venit ".
2SAM|18|28|Clamans autem Achimaas dixit ad regem: " Pax! ". Et adorans regem pronus in terram ait: " Benedictus Dominus Deus tuus, qui conclusit homines, qui levaverunt manus suas contra dominum meum regem! ".
2SAM|18|29|Et ait rex: " Estne pax puero Absalom? ". Dixitque Achimaas: " Vidi tumultum magnum, cum mitteret Ioab servum regis et me servum tuum, sed nescio quid fuerit ".
2SAM|18|30|Ad quem rex: " Recede, ait, et sta illic ". Cumque ille recessisset et staret,
2SAM|18|31|apparuit Aethiops et veniens ait: " Bonum apporto nuntium, domine mi rex; iudicavit enim pro te Dominus hodie salvans te de manu omnium, qui surrexerunt contra te ".
2SAM|18|32|Dixit autem rex ad Aethiopem: " Estne pax puero Absalom? ". Cui respondens Aethiops: " Fiant, inquit, sicut puer inimici domini mei regis et universi, qui consurrexerunt adversus eum in malum! ".
2SAM|19|1|Contremuit itaque rex et ascendit cenaculum portae et flevit. Et sic loquebatur vadens: " Fili mi Absalom, fili mi, fili mi Absalom! Quis mihi tribuat, ut ego moriar pro te? Absalom fili mi, fili mi! ".
2SAM|19|2|Nuntiatum est autem Ioab quod rex fleret et lugeret filium suum.
2SAM|19|3|Et versa est victoria in die illa in luctum omni populo; audivit enim populus in die illa dici: " Dolet rex super filio suo ".
2SAM|19|4|Et furtim ingressus est populus in die illa civitatem, quomodo reverti solet populus confusus, cum fugit de proelio.
2SAM|19|5|Porro rex operuit vultum suum et clamabat voce magna: " Fili mi Absalom, Absalom fili mi, fili mi! ".
2SAM|19|6|Ingressus ergo Ioab ad regem in domo dixit: " Confudisti hodie vultus omnium servorum tuorum, qui salvam fecerunt animam tuam hodie et animam filiorum tuorum et filiarum tuarum et animam uxorum tuarum et animam concubinarum tuarum.
2SAM|19|7|Diligis odientes te et odio habes diligentes te. Ostendisti hodie quia non curas de ducibus tuis et de servis tuis; et vere cognovi modo quia, si Absalom viveret, et nos omnes occubuissemus, tunc placeret tibi.
2SAM|19|8|Nunc igitur surge et procede et loquere ad cor servorum tuorum; iuro enim tibi per Dominum quod si non exieris, ne unus quidem remansurus sit tecum nocte hac, et peius erit hoc tibi quam omnia mala, quae venerunt super te ab adulescentia tua usque in praesens ".
2SAM|19|9|Surrexit ergo rex et sedit in porta, et omni populo nuntiatum est quod rex sederet in porta; venitque universa multitudo coram rege.Israel autem fugerat in tabernacula sua.
2SAM|19|10|Omnis quoque populus certabat in cunctis tribubus Israel dicens: " Rex liberavit nos de manu inimicorum nostrorum, ipse salvavit nos de manu Philisthinorum; et nunc fugit de terra ab Absalom.
2SAM|19|11|Absalom autem, quem unximus super nos, mortuus est in bello. Quare nunc siletis et non reducitis regem? ".
2SAM|19|12|Sermo autem omnis Israel pervenerat ad regem in domo eius. Tunc rex David misit ad Sadoc et Abiathar sacerdotes dicens: " Loquimini ad maiores natu Iudae dicentes: Cur estis novissimi ad reducendum regem in domum suam?
2SAM|19|13|Fratres mei vos, os meum et caro mea vos; quare novissimi reducitis regem?
2SAM|19|14|Et Amasae dicite: Nonne os meum es et caro mea? Haec faciat mihi Deus et haec addat, si non magister militiae fueris coram me omni tempore pro Ioab! ".
2SAM|19|15|Et inclinavit cor omnium virorum Iudae quasi viri unius; miseruntque ad regem dicentes: " Revertere tu et omnes servi tui ".
2SAM|19|16|Et reversus est rex et venit usque ad Iordanem; et Iuda venit in Galgala, ut occurreret regi et traduceret eum Iordanem.
2SAM|19|17|Festinavit autem Semei filius Gera Beniaminita de Bahurim et descendit cum viris Iudae in occursum regis David;
2SAM|19|18|mille viri de Beniamin et Siba puer de domo Saul et quindecim filii eius ac viginti servi erant cum eo. Irruperant autem Iordanem iam ante regem
2SAM|19|19|et transierant vada, ut traducerent domum regis et facerent iuxta placitum eius. Semei autem filius Gera prostratus coram rege, cum transiturus esset Iordanem,
2SAM|19|20|dixit ad eum: " Ne reputes mihi, domine mi, iniquitatem neque memineris iniuriam servi tui in die, qua egressus es, domine mi rex, de Ierusalem; neque ponas, rex, in corde tuo.
2SAM|19|21|Agnosco enim servus tuus peccatum meum et idcirco hodie primus veni de omni domo Ioseph descendique in occursum domini mei regis ".
2SAM|19|22|Respondens vero Abisai filius Sarviae dixit: " Numquid non occidetur Semei, pro hoc quia maledixit christo Domini? ".
2SAM|19|23|Et ait David: " Quid mihi et vobis, filii Sarviae, quia efficimini mihi hodie in satan? Ergone hodie interficietur vir in Israel? An ignoro hodie me factum regem super Israel? ".
2SAM|19|24|Et ait rex Semei: " Non morieris! ". Iuravitque ei.
2SAM|19|25|Meribbaal quoque filius Saul descendit in occursum regis; non laverat pedes nec circumcidit ungues nec totonderat barbam vestesque suas non laverat a die, qua egressus fuerat rex, usque ad diem reversionis eius in pace.
2SAM|19|26|Cumque de Ierusalem occurrisset regi, dixit ei rex: " Quare non venisti mecum, Meribbaal? ".
2SAM|19|27|Qui respondens ait: " Domine mi rex, servus meus decepit me! Nam dixeram ei ego famulus tuus: Sternere faciam mihi asinum et ascendens abibo cum rege; claudus enim sum servus tuus.
2SAM|19|28|Insuper et fraudulenter accusavit me servum tuum ad te dominum meum regem. Tu autem, domine mi rex, sicut angelus Dei es; fac, quod placitum est tibi.
2SAM|19|29|Neque enim fuit domus patris mei nisi morti obnoxia domino meo regi; tu autem posuisti me servum tuum inter convivas mensae tuae. Quid ultra igitur habeo iustitiae, ut vociferer ad regem? ".
2SAM|19|30|Ait ergo ei rex: " Quid ultra loqueris? Dixi: Tu et Siba dividite possessiones ".
2SAM|19|31|Responditque Meribbaal regi: " Etiam cuncta accipiat, postquam reversus est dominus meus rex pacifice in domum suam! ".
2SAM|19|32|Berzellai quoque Galaadites descenderat de Rogelim et traduxit regem Iordanem, ut dimitteret eum ad Iordanem.
2SAM|19|33|Erat autem Berzellai Galaadites senex valde, id est octogenarius; et ipse praebuerat alimenta regi, cum moraretur in Mahanaim; erat quippe vir dives nimis.
2SAM|19|34|Dixit itaque rex ad Berzellai: " Veni mecum et praebebo tibi alimenta apud me in Ierusalem ".
2SAM|19|35|Et ait Berzellai ad regem: " Quot sunt dies annorum vitae meae, ut ascendam cum rege Ierusalem?
2SAM|19|36|Octogenarius sum hodie; numquid vigent sensus mei ad discernendum suave aut amarum? Aut delectare potest servum tuum cibus et potus? Vel audire ultra possum vocem cantorum atque cantricum? Quare servus tuus esset ultra oneri domino meo regi?
2SAM|19|37|Paululum procedam famulus tuus ab Iordane tecum. Et cur dabit rex mihi hanc vicissitudinem?
2SAM|19|38|Sed obsecro, ut revertar servus tuus et moriar in civitate mea iuxta sepulcrum patris mei et matris meae. Sed ecce servus tuus Chamaam; ipse vadat tecum, domine mi rex, et fac ei, quod tibi bonum videtur ".
2SAM|19|39|Dixitque rex: " Mecum transeat Chamaam, et ego faciam ei, quidquid tibi placuerit; et omne, quod petieris a me, impetrabis ".
2SAM|19|40|Cumque transisset universus populus et rex Iordanem, osculatus est rex Berzellai et benedixit ei; et ille reversus est in locum suum.
2SAM|19|41|Transivit ergo rex in Galgala, et Chamaam cum eo. Omnis autem populus Iudae traduxerat regem, et etiam media pars populi Israel.
2SAM|19|42|Et ecce omnes viri Israel concurrentes ad regem dixerunt ei: " Quare te furati sunt fratres nostri viri Iudae et traduxerunt regem et domum eius Iordanem omnesque viros David cum eo? ".
2SAM|19|43|Et respondit omnis vir Iudae ad virum Israel: " Quia propior mihi est rex. Cur irasceris super hac re? Numquid comedimus aliquid ex rege, aut munera nobis data sunt? ".
2SAM|19|44|Et respondit vir Israel ad virum Iudae et ait: " Decem partes mihi sunt in rege et ideo etiam in David. Ego sum potior te; cur contempsisti me? Et non ego prior locutus sum, ut reducerem regem meum? ". Durius autem responderunt viri Iudae viris Israel.
2SAM|20|1|Accidit quoque, ut ibi esset vir Belial nomine Seba filius Bochri Beniaminita; et cecinit bucina et ait: Non est nobis pars in David,neque hereditas in filio Isai!Vir Israel, in tabernacula tua! ".
2SAM|20|2|Et separatus est omnis vir Israel a David secutusque est Seba filium Bochri; viri autem Iudae adhaeserunt regi suo a Iordane usque Ierusalem.
2SAM|20|3|Cumque venisset rex in domum suam Ierusalem, tulit decem mulieres concubinas, quas dereliquerat ad custodiendam domum, et tradidit eas in custodiam alimenta eis praebens. Et non est ingressus ad eas, sed erant clausae usque ad diem mortis suae in viduitate viventes.
2SAM|20|4|Dixit autem rex Amasae: " Convoca mihi omnes viros Iudae in diem tertium et tu adesto praesens ".
2SAM|20|5|Abiit ergo Amasa, ut convocaret Iudam; et moratus est ultra tempus, quod ei constituerat.
2SAM|20|6|Ait autem David ad Abisai: " Nunc magis afflicturus est nos Seba filius Bochri quam Absalom; tolle igitur servos domini tui et persequere eum, ne inveniat civitates munitas et effugiat nos ".
2SAM|20|7|Egressi sunt ergo cum eo viri Ioab, Cherethi quoque et Phelethi et omnes fortissimi; exierunt de Ierusalem ad persequendum Seba filium Bochri.
2SAM|20|8|Cumque illi essent iuxta lapidem grandem, qui est in Gabaon, Amasa venerat ante eos. Porro Ioab accinctus erat habitu suo, et in cingulo super lumbos gladius absconditus erat, qui levi motu ex vagina in manum suam cecidit.
2SAM|20|9|Dixitque Ioab ad Amasam: " Estne pax tibi, mi frater? ". Et tenuit manu dextera mentum Amasae, ut oscularetur eum.
2SAM|20|10|Porro Amasa non observavit gladium in manu Ioab, qui percussit eum in inguine et effudit intestina eius in terram, nec secundum vulnus apposuit; et mortuus est. Ioab autem et Abisai frater eius persecuti sunt Seba filium Bochri.
2SAM|20|11|Interea quidam de pueris Ioab stetit iuxta cadaver Amasae et dixit: " Qui esse vult cum Ioab et pro David, sequatur Ioab! ".
2SAM|20|12|Amasa autem conspersus sanguine iacebat in media via. Vidit hoc vir quod subsisteret omnis populus ad videndum eum; et amovit Amasam de via in agrum operuitque eum vestimento, cum videret quod omnes transeuntes propter eum subsisterent.
2SAM|20|13|Amoto igitur illo de via, transibat omnis vir sequens Ioab ad persequendum Seba filium Bochri.
2SAM|20|14|Porro ille transierat per omnes tribus Israel usque in Abelbethmaacha; omnesque Bochritae congregati sunt et ingressi sunt etiam post eum.
2SAM|20|15|Venerunt itaque et oppugnabant eum in Abelbethmaacha et fuderunt contra civitatem aggerem, qui stetit contra antemurale; et omnis populus, qui erat cum Ioab, moliebatur destruere muros.
2SAM|20|16|Et exclamavit mulier sapiens de civitate: " Audite, audite! Dicite Ioab: "Appropinqua huc, et loquar tecum" ".
2SAM|20|17|Qui cum accessisset ad eam, ait illi: " Tu es Ioab? ". Et ille respondit: " Ego ". Ad quem sic locuta est: " Audi sermones ancillae tuae. Qui respondit: " Audio ".
2SAM|20|18|Rursumque illa: " Sermo, inquit, dicebatur in vetere proverbio: Interrogent in Abel, et sic perficient rem".
2SAM|20|19|Ego pacifica fidelium Israel, et tu quaeris subruere civitatem et evertere matrem in Israel. Quare praecipitas hereditatem Domini? ".
2SAM|20|20|Respondensque Ioab ait: " Absit, absit hoc a me; non praecipito neque demolior.
2SAM|20|21|Non se sic habet res, sed homo de monte Ephraim, Seba filius Bochri cognomine, levavit manum suam contra regem David; tradite illum solum, et recedam a civitate". Et ait mulier ad Ioab: " Ecce, caput eius mittetur ad te per murum ".
2SAM|20|22|Ingressa est ergo ad omnem populum et locuta est eis sapienter. Qui abscissum caput Seba filii Bochri proiecerunt ad Ioab. Et ille cecinit tuba, et recesserunt ab urbe unusquisque in tabernacula sua. Ioab autem reversus est Ierusalem ad regem.
2SAM|20|23|Erat ergo Ioab super omnem exercitum Israel; Banaias autem filius Ioiadae super Cherethaeos et Phelethaeos;
2SAM|20|24|Adoniram vero super onera; porro Iosaphat filius Ahilud a commentariis.
2SAM|20|25|Siva autem scriba, Sadoc vero et Abiathar sacerdotes;
2SAM|20|26|Hira quoque Iairites erat sacerdos David.
2SAM|21|1|Facta est fames in diebus David tribus annis iugiter. Et consuluit David oraculum Domini, dixitque Dominus: " Super Saul et super domum eius est sanguis, quia occidit Gabaonitas ".
2SAM|21|2|Vocatis ergo Gabaonitis, rex dixit ad eos - porro Gabaonitae non sunt de filiis Israel, sed reliquiae Amorraeorum; filii quippe Israel iuraverant eis, sed voluit Saul percutere eos zelo suo pro filiis Israel et Iudae -;
2SAM|21|3|dixit ergo David ad Gabaonitas: " Quid faciam vobis? Et quod erit vestri piaculum, ut benedicatis hereditati Domini? ".
2SAM|21|4|Dixeruntque ei Gabaonitae: " Non est nobis super argento et auro quaestio contra Saul et contra domum eius; neque nobis licet interficere hominem de Israel ". Ad quos ait: " Quod ergo dixeritis, faciam vobis ".
2SAM|21|5|Qui dixerunt regi: " De filiis viri, qui attrivit nos et cogitavit delere nos ita ut ne unus quidem nostrum residuus esset in cunctis finibus Israel,
2SAM|21|6|dentur nobis septem viri, et suspendamus eos in patibulis Domino in Gabaon in monte Domini ". Et ait rex: " Ego dabo ".
2SAM|21|7|Pepercitque rex Meribbaal filio Ionathan filii Saul propter iusiurandum Domini, quod fuerat inter David et inter Ionathan filium Saul.
2SAM|21|8|Tulit itaque rex duos filios Respha filiae Aia, quos peperit Saul, Armoni et Meribbaal, et quinque filios Merob filiae Saul, quos genuerat Hadrieli filio Berzellai, qui fuit de Molathi,
2SAM|21|9|et dedit eos in manu Gabaonitarum, qui suspenderunt illos in monte coram Domino. Et ceciderunt hi septem simul, occisi in diebus messis primis, incipiente messione hordei.
2SAM|21|10|Tollens autem Respha filia Aia cilicium substravit sibi super petram ab initio messis, donec stillaret aqua super eos de caelo, et non dimisit aves caeli considere super eos per diem neque bestias campi per noctem.
2SAM|21|11|Et nuntiata sunt David, quae fecerat Respha filia Aia concubina Saul.
2SAM|21|12|Et abiit David et tulit ossa Saul et ossa Ionathan filii eius a civibus Iabes Galaad, qui furati fuerant ea de platea Bethsan, in qua suspenderant eos Philisthim, cum interfecissent Saul in Gelboe,
2SAM|21|13|et asportavit inde ossa Saul et ossa Ionathan filii eius; et colligentes ossa eorum, qui suspensi fuerant,
2SAM|21|14|sepelierunt ea cum ossibus Saul et Ionathan filii eius in terra Beniamin in Sela, in sepulcro Cis patris eius. Feceruntque omnia, quae praeceperat rex; et repropitiatus est Deus terrae post haec.
2SAM|21|15|Factum est autem rursum proelium Philisthinorum adversum Israel, et descendit David et servi eius cum eo, et pugnabant contra Philisthim, et fatigatus est David.
2SAM|21|16|Iesbibenob, qui fuit de genere Rapha - ferrum hastae trecentos siclos appendebat - et accinctus erat ense novo, nisus est percutere David;
2SAM|21|17|praesidioque ei fuit Abisai filius Sarviae et percussum Philisthaeum interfecit. Tunc iuraverunt viri David dicentes: " Iam non egredieris nobiscum in bellum, ne exstinguas lucernam Israel ".
2SAM|21|18|Fuitque rursum bellum in Gob contra Philisthaeos; tunc percussit Sobbochai de Husa Saph de stirpe Rapha.
2SAM|21|19|Et fuit iterum bellum in Gob contra Philisthaeos, in quo percussit Elchanan filius Iair Bethlehemites Goliath Getthaeum, cuius hastile hastae erat quasi liciatorium texentium.
2SAM|21|20|Et adhuc fuit bellum in Geth, in quo vir excelsus, qui senos in manibus pedibusque habebat digitos, id est viginti et quattuor, et is quoque erat de origine Rapha,
2SAM|21|21|exprobravit Israel; percussit autem eum Ionathan filius Samma fratris David.
2SAM|21|22|Hi quattuor erant de genere Rapha ex Geth et ceciderunt per manum David et servorum eius.
2SAM|22|1|Locutus est autem David Domino verba carminis huius in die, qua liberavit eum Dominus de manu omnium inimicorum suorum et de manu Saul,
2SAM|22|2|et ait: Dominus petra mea et arx mea et salvator meus;
2SAM|22|3|Deus meus, rupes mea, in quam confugiam,scutum meum et cornu salutis meae!Munimentum meum et refugium meum.Salvator meus, de violentia liberabis me.
2SAM|22|4|Laudabilem invocabo Dominumet ab inimicis meis salvus ero.
2SAM|22|5|Quia circumdederunt me fluctus mortis,torrentes Belial terruerunt me;
2SAM|22|6|praeoccupaverunt me laquei mortis.
2SAM|22|7|In tribulatione mea invocavi Dominumet ad Deum meum clamavi;et exaudivit de templo suo vocem meam,et clamor meus venit ad aures eius.
2SAM|22|8|Commota est et contremuit terra;fundamenta caelorum concussa suntet conquassata, quoniam iratus est.
2SAM|22|9|Ascendit fumus de naribus eius,et ignis de ore eius vorabat;carbones incensi sunt ab eo.
2SAM|22|10|Et inclinavit caelos et descendit,et caligo sub pedibus eius.
2SAM|22|11|Et ascendit super cherub et volavitet devolavit super pennas venti.
2SAM|22|12|Posuit tenebras in circuitu suo tabernaculum suum,tenebrosas aquas, nubes densissimas.
2SAM|22|13|Prae fulgore in conspectu eiusincensi sunt carbones ignis.
2SAM|22|14|Intonuit de caelo Dominus,et Excelsus dedit vocem suam.
2SAM|22|15|Misit sagittas et dissipavit eos,fulguravit fulmina et conturbavit eos.
2SAM|22|16|Et apparuerunt effusiones maris,et revelata sunt fundamenta orbisab increpatione Domini,ab inspiratione spiritus furoris eius.
2SAM|22|17|Misit de excelso et assumpsit me,traxit me de aquis multis;
2SAM|22|18|liberavit me ab inimico meo potentissimo,ab his, qui oderant me, qui robustiores me erant.
2SAM|22|19|Praevenerunt me in die afflictionis meae,et factus est Dominus firmamentum meum;
2SAM|22|20|et eduxit me in latitudinem,liberavit me, quia complacui ei.
2SAM|22|21|Retribuit mihi Dominus secundum iustitiam meamet secundum munditiam manuum mearum reddit mihi,
2SAM|22|22|quia custodivi vias Dominiet non egi impie a Deo meo.
2SAM|22|23|Omnia enim iudicia eius in conspectu meo,et a praeceptis eius non recessi;
2SAM|22|24|et fui immaculatus cum eoet custodivi me ab iniquitate mea.
2SAM|22|25|Et retribuet mihi Dominus secundum iustitiam meamet secundum munditiam meam in conspectu oculorum suorum.
2SAM|22|26|Cum sancto sanctus eriset cum viro innocente innocens eris;
2SAM|22|27|cum electo electus eriset cum perverso callidus eris.
2SAM|22|28|Et populum pauperem salvum facieset oculos superborum humiliabis,
2SAM|22|29|quia tu lucerna mea, Domine,et Deus meus illuminat tenebras meas.
2SAM|22|30|In te enim aggrediar hostium turmas,in Deo meo transiliam murum.
2SAM|22|31|Deus, immaculata via eius,eloquium Domini igne examinatum;scutum est omnium sperantium in se.
2SAM|22|32|Quoniam quis est Deus praeter Dominum?Et quae rupes praeter Deum nostrum?
2SAM|22|33|Deus, qui accinxit me fortitudineet complanavit perfectam viam meam,
2SAM|22|34|coaequans pedes meos cerviset super excelsa statuens me;
2SAM|22|35|docens manus meas ad proelium,et tendunt arcum aereum brachia mea.
2SAM|22|36|Dedisti mihi clipeum salutis tuae,et exauditio tua magnificavit me.
2SAM|22|37|Dilatasti gressus meos subtus me,et non sunt infirmati tali mei.
2SAM|22|38|Persequebar inimicos meos et conterebamet non convertebar, donec consumerem eos.
2SAM|22|39|Consumpsi eos et confregi, ut non consurgerent:ceciderunt sub pedibus meis.
2SAM|22|40|Accinxisti me fortitudine ad proelium,incurvasti insurgentes in me subtus me.
2SAM|22|41|Inimicos meos dedisti mihi dorsum,odientes me, et disperdidi eos.
2SAM|22|42|Clamaverunt, et non erat qui salvaret,ad Dominum, et non exaudivit eos.
2SAM|22|43|Contrivi eos ut pulverem terrae,quasi lutum platearum comminui eos.
2SAM|22|44|Salvasti me a contradictionibus populi mei,constituisti me in caput gentium.Populus, quem ignorabam, servit mihi,
2SAM|22|45|filii alieni blandiuntur mihi,auditu auris oboediunt mihi.
2SAM|22|46|Filii alieni defluuntet contremiscunt ex arcibus suis.
2SAM|22|47|Vivit Dominus, et benedicta petra mea,et exaltetur Deus, petra salutis meae.
2SAM|22|48|Deus, qui das vindictas mihiet deicis populos sub me.
2SAM|22|49|Qui educis me ab inimicis meiset ab insurgentibus in me elevas me;a viro iniquo liberas me.
2SAM|22|50|Propterea confitebor tibi, Domine, in gentibus,et nomini tuo cantabo:
2SAM|22|51|Magnificat salutes regis suiet facit misericordiam christo suo Davidet semini eius in sempiternum ".
2SAM|23|1|Haec autem sunt verba David novissima: Dixit David filius Isai,dixit vir constitutus in alto,christus Dei Iacob,suavis psalta Israel.
2SAM|23|2|Spiritus Domini locutus est per me, et sermo eius super linguam meam.
2SAM|23|3|Locutus est Deus Israel,mihi dixit Petra Israel:Dominator hominum iustus,dominator in timore Dei
2SAM|23|4|est sicut lux aurorae, oriente sole,mane absque nubibus;de splendore post pluviamherba oritur de terra".
2SAM|23|5|Nonne sic est domus mea cum Deo?Quia pactum aeternum statuit mihi,dispositum in omnibus atque munitum.Cunctam enim salutem meam et omne desiderabilenonne faciet germinare?
2SAM|23|6|Praevaricatores autemquasi spinae abiectae universi,quae non tolluntur manibus;
2SAM|23|7|et si quis tangere voluerit eas,armabitur ferro et ligno lanceato,igneque succensae comburentur ".
2SAM|23|8|Haec nomina fortium David:Iesbaal Hachamonites, princeps inter tres, ipse levavit hastam suam super octingentos, quos interfecit impetu uno.
2SAM|23|9|Post hunc Eleazar filius Dodo Ahohites, inter tres fortes. Qui erat cum David in Aphesdommim, quando Philisthim congregati sunt illuc in proelium.
2SAM|23|10|Cumque ascendissent viri Israel, ipse stetit et percussit Philisthaeos, donec deficeret manus eius et obrigesceret cum gladio; fecitque Dominus salutem magnam in die illa, et populus reversus est tantum ad spolia detrahenda.
2SAM|23|11|Et post hunc Samma filius Age Ararites. Et congregati sunt Philisthim in Lehi; erat quippe ibi ager lente plenus. Cumque fugisset populus a facie Philisthim,
2SAM|23|12|stetit ille in medio agri et tuitus est eum percussitque Philisthaeos, et fecit Dominus salutem magnam.
2SAM|23|13|Et descenderunt tres de triginta et venerunt tempore messis ad David in speluncam Odollam; castra autem Philisthinorum erant posita in valle Raphaim.
2SAM|23|14|Et David erat tunc in praesidio; porro statio Philisthinorum tunc erat in Bethlehem.
2SAM|23|15|Desideravit igitur David et ait: " O si quis mihi daret potum aquae de cisterna, quae est in Bethlehem iuxta portam! ".
2SAM|23|16|Irruperunt ergo tres fortes castra Philisthinorum et hauserunt aquam de cisterna Bethlehem, quae erat iuxta portam, et attulerunt ad David. At ille noluit bibere, sed libavit illam Domino
2SAM|23|17|dicens: " Propitius mihi sit Dominus, ne faciam hoc. Num sanguinem hominum istorum, qui profecti sunt in animarum periculo, bibam? ". Noluit ergo bibere. Haec fecerunt tres robustissimi.
2SAM|23|18|Abisai autem frater Ioab filius Sarviae princeps erat de triginta. Ipse est qui elevavit hastam suam contra trecentos, quos interfecit. Nominatus in triginta
2SAM|23|19|et inter triginta nobilior eratque eorum princeps; sed usque ad tres primos non pervenerat.
2SAM|23|20|Et Banaias filius Ioiadae vir fortissimus magnorum operum de Cabseel. Ipse percussit duos filios Ariel de Moab, et ipse descendit et percussit leonem in media cisterna in diebus nivis.
2SAM|23|21|Ipse quoque interfecit virum Aegyptium, virum procerae staturae habentem in manu hastam; itaque cum descendisset ad eum cum baculo, vi extorsit hastam de manu Aegyptii et interfecit eum hasta sua.
2SAM|23|22|Haec fecit Banaias filius Ioiadae, et ipse nominatus inter triginta fortissimos.
2SAM|23|23|Erat autem nobilior inter triginta; verumtamen usque ad tres non pervenerat. Fecitque eum David sibi caput satellitum suorum.
2SAM|23|24|Asael frater Ioab erat inter triginta. Elchanan filius Dodo de Bethlehem,
2SAM|23|25|Samma de Harod, Elica de Harod,
2SAM|23|26|Heles de Phalti, Hira filius Acces de Thecua,
2SAM|23|27|Abiezer de Anathoth, Sobbochai de Husa,
2SAM|23|28|Selmon Ahohites, Maharai Netophathites,
2SAM|23|29|Heled filius Baana Netophathites, Ithai filius Ribai de Gabaa filiorum Beniamin,
2SAM|23|30|Banaia Pharathonites, Heddai de torrentibus Gaas,
2SAM|23|31|Abibaal Arbathites, Azmaveth de Bahurim,
2SAM|23|32|Eliaba de Saalbon, Iasen de Gun,
2SAM|23|33|Ionathan filius Samma de Arar, Ahiam filius Sarar Ararites.
2SAM|23|34|Eliphalet filius Aasbai Maachathitae, Eliam filius Achitophel Gilonites,
2SAM|23|35|Hesro de Carmel, Pharai de Arab,
2SAM|23|36|Igal filius Nathan de Soba, Bani de Gad,
2SAM|23|37|Selec de Ammon, Naharai Berothites armiger Ioab filii Sarviae,
2SAM|23|38|Hira Iethrites, Gareb et ipse Iethrites,
2SAM|23|39|Urias Hetthaeus.Omnes triginta septem.
2SAM|24|1|Et addidit furor Domini ira sci contra Israel; commovit que David contra eos dicens: " Vade, numera Israel et Iudam ".
2SAM|24|2|Dixitque rex ad Ioab et ad principes exercitus sui, qui erant cum eo: " Perambula omnes tribus Israel a Dan usque Bersabee, et numerate populum, ut sciam numerum eius ".
2SAM|24|3|Dixitque Ioab regi: " Adaugeat Dominus Deus tuus ad populum, quantus nunc est, centuplum in conspectu domini mei regis! Sed quid sibi dominus meus rex vult in re huiuscemodi? ".
2SAM|24|4|Praevaluit autem sermo regis contra Ioab et principes exercitus; egressusque est Ioab et principes militum a facie regis, ut numerarent populum Israel.
2SAM|24|5|Cumque pertransissent Iordanem, inceperunt ab Aroer et ab urbe, quae est in media valle, transeuntes ad Gaditas et ad Iazer.
2SAM|24|6|Et pervenerunt in Galaad et in terram Hetthaeorum in Cades et venerunt in Dan. Et a Dan converterunt se ad Sidonem
2SAM|24|7|et pervenerunt ad arcem Tyri et omnes urbes Hevaei et Chananaei exieruntque ad Nageb Iudae in Bersabee.
2SAM|24|8|Et, lustrata universa terra, affuerunt post novem menses et viginti dies in Ierusalem.
2SAM|24|9|Dedit ergo Ioab numerum descriptionis populi regi; et inventa sunt de Israel octingenta milia virorum fortium, qui educerent gladium, et de Iuda quingenta milia pugnatorum.
2SAM|24|10|Percussit autem cor David eum, postquam numeratus est populus, et dixit David ad Dominum: " Peccavi valde in hoc facto; nunc vero precor, Domine, ut transferas iniquitatem servi tui, quia stulte egi nimis ".
2SAM|24|11|Surrexit itaque David mane, et sermo Domini factus est ad Gad propheten, videntem David, dicens:
2SAM|24|12|" Vade et loquere ad David: Haec dicit Dominus: Trium tibi datur optio; elige unum, quod volueris ex his, ut faciam tibi ".
2SAM|24|13|Cumque venisset Gad ad David, nuntiavit ei dicens: " Aut tribus annis veniet tibi fames in terra tua, aut tribus mensibus fugies adversarios tuos, et illi te persequentur, aut certe tribus diebus erit pestilentia in terra tua. Nunc ergo delibera et vide quem respondeam ei, qui me misit, sermonem ".
2SAM|24|14|Dixit autem David ad Gad: " Artor nimis; sed melius est, ut incidamus in manu Domini - multae enim misericordiae eius sunt - quam in manu hominum! ".
2SAM|24|15|Et elegit sibi David pestilentiam; et erant dies messis tritici. Immisitque Dominus pestilentiam in Israel de mane usque ad tempus constitutum, et mortui sunt ex populo a Dan usque Bersabee septuaginta milia virorum.
2SAM|24|16|Cumque extendisset manum suam angelus super Ierusalem, ut disperderet eam, misertus est Dominus super afflictione et ait angelo percutienti populum: " Sufficit; nunc contine manum tuam! ".Erat autem angelus Domini iuxta aream Areuna Iebusaei.
2SAM|24|17|Dixitque David ad Dominum, cum vidisset angelum caedentem populum: " Ego sum qui peccavi, ego inique egi; isti, qui oves sunt, quid fecerunt? Vertatur, obsecro, manus tua contra me et contra domum patris mei ".
2SAM|24|18|Venit autem Gad ad David in die illa et dixit ei: " Ascende, constitue Domino altare in area Areuna Iebusaei ".
2SAM|24|19|Et ascendit David iuxta sermonem Gad, quem praeceperat ei Dominus.
2SAM|24|20|Conspiciensque Areuna animadvertit regem et servos eius transire ad se
2SAM|24|21|et egressus adoravit regem prono vultu in terra et ait: " Quid causae est, ut veniat dominus meus rex ad servum suum? ". Cui David ait: " Ut emam a te aream et aedificem altare Domino, et cesset interfectio, quae grassatur in populo ".
2SAM|24|22|Et ait Areuna ad David: " Accipiat et offerat dominus meus rex, sicut ei placet. Ecce boves in holocaustum et plaustrum et iuga boum in usum lignorum.
2SAM|24|23|Omnia dat Areuna, o rex, regi ". Dixitque Areuna ad regem: " Dominus Deus tuus suscipiat votum tuum! ".
2SAM|24|24|Cui respondens rex ait: " Nequaquam; sed emam pretio a te et non offeram Domino Deo meo holocausta gratuita ". Emit ergo David aream et boves argenti siclis quinquaginta.
2SAM|24|25|Et aedificavit ibi David altare Domino et obtulit holocausta et pacifica.Et repropitiatus est Dominus terrae, et cohibita est plaga ab Israel.
