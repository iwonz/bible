2PET|1|1|Simeon Peter, a servant and apostle of Jesus Christ, To those who have obtained a faith of equal standing with ours by the righteousness of our God and Savior Jesus Christ:
2PET|1|2|May grace and peace be multiplied to you in the knowledge of God and of Jesus our Lord.
2PET|1|3|His divine power has granted to us all things that pertain to life and godliness, through the knowledge of him who called us to his own glory and excellence,
2PET|1|4|by which he has granted to us his precious and very great promises, so that through them you may become partakers of the divine nature, having escaped from the corruption that is in the world because of sinful desire.
2PET|1|5|For this very reason, make every effort to supplement your faith with virtue, and virtue with knowledge,
2PET|1|6|and knowledge with self-control, and self-control with steadfastness, and steadfastness with godliness,
2PET|1|7|and godliness with brotherly affection, and brotherly affection with love.
2PET|1|8|For if these qualities are yours and are increasing, they keep you from being ineffective or unfruitful in the knowledge of our Lord Jesus Christ.
2PET|1|9|For whoever lacks these qualities is so nearsighted that he is blind, having forgotten that he was cleansed from his former sins.
2PET|1|10|Therefore, brothers, be all the more diligent to make your calling and election sure, for if you practice these qualities you will never fall.
2PET|1|11|For in this way there will be richly provided for you an entrance into the eternal kingdom of our Lord and Savior Jesus Christ.
2PET|1|12|Therefore I intend always to remind you of these qualities, though you know them and are established in the truth that you have.
2PET|1|13|I think it right, as long as I am in this body, to stir you up by way of reminder,
2PET|1|14|since I know that the putting off of my body will be soon, as our Lord Jesus Christ made clear to me.
2PET|1|15|And I will make every effort so that after my departure you may be able at any time to recall these things.
2PET|1|16|For we did not follow cleverly devised myths when we made known to you the power and coming of our Lord Jesus Christ, but we were eyewitnesses of his majesty.
2PET|1|17|For when he received honor and glory from God the Father, and the voice was borne to him by the Majestic Glory, "This is my beloved Son, with whom I am well pleased,"
2PET|1|18|we ourselves heard this very voice borne from heaven, for we were with him on the holy mountain.
2PET|1|19|And we have something more sure, the prophetic word, to which you will do well to pay attention as to a lamp shining in a dark place, until the day dawns and the morning star rises in your hearts,
2PET|1|20|knowing this first of all, that no prophecy of Scripture comes from someone's own interpretation.
2PET|1|21|For no prophecy was ever produced by the will of man, but men spoke from God as they were carried along by the Holy Spirit.
2PET|2|1|But false prophets also arose among the people, just as there will be false teachers among you, who will secretly bring in destructive heresies, even denying the Master who bought them, bringing upon themselves swift destruction.
2PET|2|2|And many will follow their sensuality, and because of them the way of truth will be blasphemed.
2PET|2|3|And in their greed they will exploit you with false words. Their condemnation from long ago is not idle, and their destruction is not asleep.
2PET|2|4|For if God did not spare angels when they sinned, but cast them into hell and committed them to chains of gloomy darkness to be kept until the judgment;
2PET|2|5|if he did not spare the ancient world, but preserved Noah, a herald of righteousness, with seven others, when he brought a flood upon the world of the ungodly;
2PET|2|6|if by turning the cities of Sodom and Gomorrah to ashes he condemned them to extinction, making them an example of what is going to happen to the ungodly;
2PET|2|7|and if he rescued righteous Lot, greatly distressed by the sensual conduct of the wicked
2PET|2|8|(for as that righteous man lived among them day after day, he was tormenting his righteous soul over their lawless deeds that he saw and heard);
2PET|2|9|then the Lord knows how to rescue the godly from trials, and to keep the unrighteous under punishment until the day of judgment,
2PET|2|10|and especially those who indulge in the lust of defiling passion and despise authority. Bold and willful, they do not tremble as they blaspheme the glorious ones,
2PET|2|11|whereas angels, though greater in might and power, do not pronounce a blasphemous judgment against them before the Lord.
2PET|2|12|But these, like irrational animals, creatures of instinct, born to be caught and destroyed, blaspheming about matters of which they are ignorant, will also be destroyed in their destruction,
2PET|2|13|suffering wrong as the wage for their wrongdoing. They count it pleasure to revel in the daytime. They are blots and blemishes, reveling in their deceptions, while they feast with you.
2PET|2|14|They have eyes full of adultery, insatiable for sin. They entice unsteady souls. They have hearts trained in greed. Accursed children!
2PET|2|15|Forsaking the right way, they have gone astray. They have followed the way of Balaam, the son of Beor, who loved gain from wrongdoing,
2PET|2|16|but was rebuked for his own transgression; a speechless donkey spoke with human voice and restrained the prophet's madness.
2PET|2|17|These are waterless springs and mists driven by a storm. For them the gloom of utter darkness has been reserved.
2PET|2|18|For, speaking loud boasts of folly, they entice by sensual passions of the flesh those who are barely escaping from those who live in error.
2PET|2|19|They promise them freedom, but they themselves are slaves of corruption. For whatever overcomes a person, to that he is enslaved.
2PET|2|20|For if, after they have escaped the defilements of the world through the knowledge of our Lord and Savior Jesus Christ, they are again entangled in them and overcome, the last state has become worse for them than the first.
2PET|2|21|For it would have been better for them never to have known the way of righteousness than after knowing it to turn back from the holy commandment delivered to them.
2PET|2|22|What the true proverb says has happened to them: "The dog returns to its own vomit, and the sow, after washing herself, returns to wallow in the mire."
2PET|3|1|This is now the second letter that I am writing to you, beloved. In both of them I am stirring up your sincere mind by way of reminder,
2PET|3|2|that you should remember the predictions of the holy prophets and the commandment of the Lord and Savior through your apostles,
2PET|3|3|knowing this first of all, that scoffers will come in the last days with scoffing, following their own sinful desires.
2PET|3|4|They will say, "Where is the promise of his coming? For ever since the fathers fell asleep, all things are continuing as they were from the beginning of creation."
2PET|3|5|For they deliberately overlook this fact, that the heavens existed long ago, and the earth was formed out of water and through water by the word of God,
2PET|3|6|and that by means of these the world that then existed was deluged with water and perished.
2PET|3|7|But by the same word the heavens and earth that now exist are stored up for fire, being kept until the day of judgment and destruction of the ungodly.
2PET|3|8|But do not overlook this one fact, beloved, that with the Lord one day is as a thousand years, and a thousand years as one day.
2PET|3|9|The Lord is not slow to fulfill his promise as some count slowness, but is patient toward you, not wishing that any should perish, but that all should reach repentance.
2PET|3|10|But the day of the Lord will come like a thief, and then the heavens will pass away with a roar, and the heavenly bodies will be burned up and dissolved, and the earth and the works that are done on it will be exposed.
2PET|3|11|Since all these things are thus to be dissolved, what sort of people ought you to be in lives of holiness and godliness,
2PET|3|12|waiting for and hastening the coming of the day of God, because of which the heavens will be set on fire and dissolved, and the heavenly bodies will melt as they burn!
2PET|3|13|But according to his promise we are waiting for new heavens and a new earth in which righteousness dwells.
2PET|3|14|Therefore, beloved, since you are waiting for these, be diligent to be found by him without spot or blemish, and at peace.
2PET|3|15|And count the patience of our Lord as salvation, just as our beloved brother Paul also wrote to you according to the wisdom given him,
2PET|3|16|as he does in all his letters when he speaks in them of these matters. There are some things in them that are hard to understand, which the ignorant and unstable twist to their own destruction, as they do the other Scriptures.
2PET|3|17|You therefore, beloved, knowing this beforehand, take care that you are not carried away with the error of lawless people and lose your own stability.
2PET|3|18|But grow in the grace and knowledge of our Lord and Savior Jesus Christ. To him be the glory both now and to the day of eternity. Amen.
