1TIM|1|1|Paulus apostolus Christi Iesu secundum imperium Dei salvatoris nostri et Christi Iesu spei nostrae
1TIM|1|2|Timotheo dilecto filio in fide gratia misericordia pax a Deo Patre et Christo Iesu Domino nostro
1TIM|1|3|sicut rogavi te ut remaneres Ephesi cum irem in Macedoniam ut denuntiares quibusdam ne aliter docerent
1TIM|1|4|neque intenderent fabulis et genealogiis interminatis quae quaestiones praestant magis quam aedificationem Dei quae est in fide
1TIM|1|5|finis autem praecepti est caritas de corde puro et conscientia bona et fide non ficta
1TIM|1|6|a quibus quidam aberrantes conversi sunt in vaniloquium
1TIM|1|7|volentes esse legis doctores non intellegentes neque quae loquuntur neque de quibus adfirmant
1TIM|1|8|scimus autem quia bona est lex si quis ea legitime utatur
1TIM|1|9|sciens hoc quia iusto lex non est posita sed iniustis et non subditis impiis et peccatoribus sceleratis et contaminatis patricidis et matricidis homicidis
1TIM|1|10|fornicariis masculorum concubitoribus plagiariis mendacibus periuris et si quid aliud sanae doctrinae adversatur
1TIM|1|11|quae est secundum evangelium gloriae beati Dei quod creditum est mihi
1TIM|1|12|gratias ago ei qui me confortavit Christo Iesu Domino nostro quia fidelem me existimavit ponens in ministerio
1TIM|1|13|qui prius fui blasphemus et persecutor et contumeliosus sed misericordiam consecutus sum quia ignorans feci in incredulitate
1TIM|1|14|superabundavit autem gratia Domini nostri cum fide et dilectione quae est in Christo Iesu
1TIM|1|15|fidelis sermo et omni acceptione dignus quia Christus Iesus venit in mundum peccatores salvos facere quorum primus ego sum
1TIM|1|16|sed ideo misericordiam consecutus sum ut in me primo ostenderet Christus Iesus omnem patientiam ad deformationem eorum qui credituri sunt illi in vitam aeternam
1TIM|1|17|regi autem saeculorum inmortali invisibili soli Deo honor et gloria in saecula saeculorum amen
1TIM|1|18|hoc praeceptum commendo tibi fili Timothee secundum praecedentes in te prophetias ut milites in illis bonam militiam
1TIM|1|19|habens fidem et bonam conscientiam quam quidam repellentes circa fidem naufragaverunt
1TIM|1|20|ex quibus est Hymeneus et Alexander quos tradidi Satanae ut discant non blasphemare
1TIM|2|1|obsecro igitur primo omnium fieri obsecrationes orationes postulationes gratiarum actiones pro omnibus hominibus
1TIM|2|2|pro regibus et omnibus qui in sublimitate sunt ut quietam et tranquillam vitam agamus in omni pietate et castitate
1TIM|2|3|hoc enim bonum est et acceptum coram salutari nostro Deo
1TIM|2|4|qui omnes homines vult salvos fieri et ad agnitionem veritatis venire
1TIM|2|5|unus enim Deus unus et mediator Dei et hominum homo Christus Iesus
1TIM|2|6|qui dedit redemptionem semet ipsum pro omnibus testimonium temporibus suis
1TIM|2|7|in quo positus sum ego praedicator et apostolus veritatem dico non mentior doctor gentium in fide et veritate
1TIM|2|8|volo ergo viros orare in omni loco levantes puras manus sine ira et disceptatione
1TIM|2|9|similiter et mulieres in habitu ornato cum verecundia et sobrietate ornantes se non in tortis crinibus aut auro aut margaritis vel veste pretiosa
1TIM|2|10|sed quod decet mulieres promittentes pietatem per opera bona
1TIM|2|11|mulier in silentio discat cum omni subiectione
1TIM|2|12|docere autem mulieri non permitto neque dominari in virum sed esse in silentio
1TIM|2|13|Adam enim primus formatus est deinde Eva
1TIM|2|14|et Adam non est seductus mulier autem seducta in praevaricatione fuit
1TIM|2|15|salvabitur autem per filiorum generationem si permanserint in fide et dilectione et sanctificatione cum sobrietate
1TIM|3|1|fidelis sermo si quis episcopatum desiderat bonum opus desiderat
1TIM|3|2|oportet ergo episcopum inreprehensibilem esse unius uxoris virum sobrium prudentem ornatum hospitalem doctorem
1TIM|3|3|non vinolentum non percussorem sed modestum non litigiosum non cupidum
1TIM|3|4|suae domui bene praepositum filios habentem subditos cum omni castitate
1TIM|3|5|si quis autem domui suae praeesse nescit quomodo ecclesiae Dei diligentiam habebit
1TIM|3|6|non neophytum ne in superbia elatus in iudicium incidat diaboli
1TIM|3|7|oportet autem illum et testimonium habere bonum ab his qui foris sunt ut non in obprobrium incidat et laqueum diaboli
1TIM|3|8|diaconos similiter pudicos non bilingues non multo vino deditos non turpe lucrum sectantes
1TIM|3|9|habentes mysterium fidei in conscientia pura
1TIM|3|10|et hii autem probentur primum et sic ministrent nullum crimen habentes
1TIM|3|11|mulieres similiter pudicas non detrahentes sobrias fideles in omnibus
1TIM|3|12|diacones sint unius uxoris viri qui filiis suis bene praesunt et suis domibus
1TIM|3|13|qui enim bene ministraverint gradum sibi bonum adquirent et multam fiduciam in fide quae est in Christo Iesu
1TIM|3|14|haec tibi scribo sperans venire ad te cito
1TIM|3|15|si autem tardavero ut scias quomodo oporteat te in domo Dei conversari quae est ecclesia Dei vivi columna et firmamentum veritatis
1TIM|3|16|et manifeste magnum est pietatis sacramentum quod manifestatum est in carne iustificatum est in spiritu apparuit angelis praedicatum est gentibus creditum est in mundo adsumptum est in gloria
1TIM|4|1|Spiritus autem manifeste dicit quia in novissimis temporibus discedent quidam a fide adtendentes spiritibus erroris et doctrinis daemoniorum
1TIM|4|2|in hypocrisi loquentium mendacium et cauteriatam habentium suam conscientiam
1TIM|4|3|prohibentium nubere abstinere a cibis quos Deus creavit ad percipiendum cum gratiarum actione fidelibus et his qui cognoverunt veritatem
1TIM|4|4|quia omnis creatura Dei bona et nihil reiciendum quod cum gratiarum actione percipitur
1TIM|4|5|sanctificatur enim per verbum Dei et orationem
1TIM|4|6|haec proponens fratribus bonus eris minister Christi Iesu enutritus verbis fidei et bonae doctrinae quam adsecutus es
1TIM|4|7|ineptas autem et aniles fabulas devita exerce te ipsum ad pietatem
1TIM|4|8|nam corporalis exercitatio ad modicum utilis est pietas autem ad omnia utilis est promissionem habens vitae quae nunc est et futurae
1TIM|4|9|fidelis sermo et omni acceptione dignus
1TIM|4|10|in hoc enim laboramus et maledicimur quia speravimus in Deum vivum qui est salvator omnium hominum maxime fidelium
1TIM|4|11|praecipe haec et doce
1TIM|4|12|nemo adulescentiam tuam contemnat sed exemplum esto fidelium in verbo in conversatione in caritate in fide in castitate
1TIM|4|13|dum venio adtende lectioni exhortationi doctrinae
1TIM|4|14|noli neglegere gratiam quae in te est quae data est tibi per prophetiam cum inpositione manuum presbyterii
1TIM|4|15|haec meditare in his esto ut profectus tuus manifestus sit omnibus
1TIM|4|16|adtende tibi et doctrinae insta in illis hoc enim faciens et te ipsum salvum facies et qui te audiunt
1TIM|5|1|seniorem ne increpaveris sed obsecra ut patrem iuvenes ut fratres
1TIM|5|2|anus ut matres iuvenculas ut sorores in omni castitate
1TIM|5|3|viduas honora quae vere viduae sunt
1TIM|5|4|si qua autem vidua filios aut nepotes habet discant primum domum suam regere et mutuam vicem reddere parentibus hoc enim acceptum est coram Deo
1TIM|5|5|quae autem vere vidua est et desolata speravit in Deum et instat obsecrationibus et orationibus nocte ac die
1TIM|5|6|nam quae in deliciis est vivens mortua est
1TIM|5|7|et hoc praecipe ut inreprehensibiles sint
1TIM|5|8|si quis autem suorum et maxime domesticorum curam non habet fidem negavit et est infideli deterior
1TIM|5|9|vidua eligatur non minus sexaginta annorum quae fuerit unius viri uxor
1TIM|5|10|in operibus bonis testimonium habens si filios educavit si hospitio recepit si sanctorum pedes lavit si tribulationem patientibus subministravit si omne opus bonum subsecuta est
1TIM|5|11|adulescentiores autem viduas devita cum enim luxuriatae fuerint in Christo nubere volunt
1TIM|5|12|habentes damnationem quia primam fidem irritam fecerunt
1TIM|5|13|simul autem et otiosae discunt circumire domos non solum otiosae sed et verbosae et curiosae loquentes quae non oportet
1TIM|5|14|volo ergo iuveniores nubere filios procreare matres familias esse nullam occasionem dare adversario maledicti gratia
1TIM|5|15|iam enim quaedam conversae sunt retro Satanan
1TIM|5|16|si qua fidelis habet viduas subministret illis et non gravetur ecclesia ut his quae vere viduae sunt sufficiat
1TIM|5|17|qui bene praesunt presbyteri duplici honore digni habeantur maxime qui laborant in verbo et doctrina
1TIM|5|18|dicit enim scriptura non infrenabis os bovi trituranti et dignus operarius mercede sua
1TIM|5|19|adversus presbyterum accusationem noli recipere nisi sub duobus et tribus testibus
1TIM|5|20|peccantes coram omnibus argue ut et ceteri timorem habeant
1TIM|5|21|testor coram Deo et Christo Iesu et electis angelis ut haec custodias sine praeiudicio nihil faciens in aliam partem declinando
1TIM|5|22|manus cito nemini inposueris neque communicaveris peccatis alienis te ipsum castum custodi
1TIM|5|23|noli adhuc aquam bibere sed vino modico utere propter stomachum tuum et frequentes tuas infirmitates
1TIM|5|24|quorundam hominum peccata manifesta sunt praecedentia ad iudicium quosdam autem et subsequuntur
1TIM|5|25|similiter et facta bona manifesta sunt et quae aliter se habent abscondi non possunt
1TIM|6|1|quicumque sunt sub iugo servi dominos suos omni honore dignos arbitrentur ne nomen Domini et doctrina blasphemetur
1TIM|6|2|qui autem fideles habent dominos non contemnant quia fratres sunt sed magis serviant quia fideles sunt et dilecti qui beneficii participes sunt haec doce et exhortare
1TIM|6|3|si quis aliter docet et non adquiescit sanis sermonibus Domini nostri Iesu Christi et ei quae secundum pietatem est doctrinae
1TIM|6|4|superbus nihil sciens sed languens circa quaestiones et pugnas verborum ex quibus oriuntur invidiae contentiones blasphemiae suspiciones malae
1TIM|6|5|conflictationes hominum mente corruptorum et qui veritate privati sunt existimantium quaestum esse pietatem
1TIM|6|6|est autem quaestus magnus pietas cum sufficientia
1TIM|6|7|nihil enim intulimus in mundum haut dubium quia nec auferre quid possumus
1TIM|6|8|habentes autem alimenta et quibus tegamur his contenti sumus
1TIM|6|9|nam qui volunt divites fieri incidunt in temptationem et laqueum et desideria multa inutilia et nociva quae mergunt homines in interitum et perditionem
1TIM|6|10|radix enim omnium malorum est cupiditas quam quidam appetentes erraverunt a fide et inseruerunt se doloribus multis
1TIM|6|11|tu autem o homo Dei haec fuge sectare vero iustitiam pietatem fidem caritatem patientiam mansuetudinem
1TIM|6|12|certa bonum certamen fidei adprehende vitam aeternam in qua vocatus es et confessus bonam confessionem coram multis testibus
1TIM|6|13|praecipio tibi coram Deo qui vivificat omnia et Christo Iesu qui testimonium reddidit sub Pontio Pilato bonam confessionem
1TIM|6|14|ut serves mandatum sine macula inreprehensibile usque in adventum Domini nostri Iesu Christi
1TIM|6|15|quem suis temporibus ostendet beatus et solus potens rex regum et Dominus dominantium
1TIM|6|16|qui solus habet inmortalitatem lucem habitans inaccessibilem quem vidit nullus hominum sed nec videre potest cui honor et imperium sempiternum amen
1TIM|6|17|divitibus huius saeculi praecipe non sublime sapere neque sperare in incerto divitiarum sed in Deo qui praestat nobis omnia abunde ad fruendum
1TIM|6|18|bene agere divites fieri in operibus bonis facile tribuere communicare
1TIM|6|19|thesaurizare sibi fundamentum bonum in futurum ut adprehendant veram vitam
1TIM|6|20|o Timothee depositum custodi devitans profanas vocum novitates et oppositiones falsi nominis scientiae
1TIM|6|21|quam quidam promittentes circa fidem exciderunt gratia tecum
