MATT|1|1|Liber generationis Iesu Christi filii David filii Abraham.
MATT|1|2|Abraham genuit Isaac, Isaac autem genuit Iacob, Iacob autem genuit Iudam et fratres eius,
MATT|1|3|Iudas autem genuit Phares et Zara de Thamar, Phares autem genuit Esrom, Esrom autem genuit Aram,
MATT|1|4|Aram autem genuit Aminadab, Aminadab autem genuit Naasson, Naasson autem genuit Salmon,
MATT|1|5|Salmon autem genuit Booz de Rahab, Booz autem genuit Obed ex Ruth, Obed autem genuit Iesse,
MATT|1|6|Iesse autem genuit David regem.David autem genuit Salomonem ex ea, quae fuit Uriae,
MATT|1|7|Salomon autem genuit Roboam, Roboam autem genuit Abiam, Abia autem genuit Asa,
MATT|1|8|Asa autem genuit Iosaphat, Iosaphat autem genuit Ioram, Ioram autem genuit Oziam,
MATT|1|9|Ozias autem genuit Ioatham, Ioatham autem genuit Achaz, Achaz autem genuit Ezechiam,
MATT|1|10|Ezechias autem genuit Manassen, Manasses autem genuit Amon, Amon autem genuit Iosiam,
MATT|1|11|Iosias autem genuit Iechoniam et fratres eius in transmigratione Babylonis.
MATT|1|12|Et post transmigrationem Babylonis Iechonias genuit Salathiel, Salathiel autem genuit Zorobabel,
MATT|1|13|Zorobabel autem genuit Abiud, Abiud autem genuit Eliachim, Eliachim autem genuit Azor,
MATT|1|14|Azor autem genuit Sadoc, Sadoc autem genuit Achim, Achim autem genuit Eliud,
MATT|1|15|Eliud autem genuit Eleazar, Eleazar autem genuit Matthan, Matthan autem genuit Iacob,
MATT|1|16|Iacob autem genuit Ioseph virum Mariae, de qua natus est Iesus, qui vocatur Christus.
MATT|1|17|Omnes ergo generationes ab Abraham usque ad David generationes quattuordecim; et a David usque ad transmigrationem Babylonis generationes quattuordecim; et a transmigratione Babylonis usque ad Christum generationes quattuordecim.
MATT|1|18|Iesu Christi autem generatio sic erat.Cum esset desponsata mater eius Maria Ioseph, antequam convenirent inventa est in utero habens de Spiritu Sancto.
MATT|1|19|Ioseph autem vir eius, cum esset iustus et nollet eam traducere, voluit occulte dimittere eam.
MATT|1|20|Haec autem eo cogitante, ecce angelus Domini in somnis apparuit ei dicens: " Ioseph fili David, noli timere accipere Mariam coniugem tuam. Quod enim in ea natum est, de Spiritu Sancto est;
MATT|1|21|pariet autem filium, et vocabis nomen eius Iesum: ipse enim salvum faciet populum suum a peccatis eorum ".
MATT|1|22|Hoc autem totum factum est, ut adimpleretur id, quod dictum est a Domino per prophetam dicentem:
MATT|1|23|" Ecce, virgo in utero habebit et pariet filium, et vocabunt nomen eius Emmanuel ", quod est interpretatum Nobiscum Deus.
MATT|1|24|Exsurgens autem Ioseph a somno fecit, sicut praecepit ei angelus Domini, et accepit coniugem suam;
MATT|1|25|et non cognoscebat eam, donec peperit filium, et vocavit nomen eius Iesum.
MATT|2|1|Cum autem natus esset Iesus in Bethlehem Iudaeae in diebus Herodis regis, ecce Magi ab oriente venerunt Hierosolymam
MATT|2|2|dicentes: " Ubi est, qui natus est, rex Iudaeorum? Vidimus enim stellam eius in oriente et venimus adorare eum ".
MATT|2|3|Audiens autem Herodes rex turbatus est et omnis Hierosolyma cum illo;
MATT|2|4|et congregans omnes principes sacerdotum et scribas populi, sciscitabatur ab eis ubi Christus nasceretur.
MATT|2|5|At illi dixerunt ei: " In Bethlehem Iudaeae. Sic enim scriptum est per prophetam:
MATT|2|6|"Et tu, Bethlehem terra Iudae,nequaquam minima es in principibus Iudae;ex te enim exiet dux,qui reget populum meum Israel" ".
MATT|2|7|Tunc Herodes, clam vocatis Magis, diligenter didicit ab eis tempus stellae, quae apparuit eis;
MATT|2|8|et mittens illos in Bethlehem dixit: " Ite et interrogate diligenter de puero; et cum inveneritis, renuntiate mihi, ut et ego veniens adorem eum.
MATT|2|9|Qui cum audissent regem, abierunt. Et ecce stella, quam viderant in oriente, antecedebat eos, usque dum veniens staret supra, ubi erat puer.
MATT|2|10|Videntes autem stellam gavisi sunt gaudio magno valde.
MATT|2|11|Et intrantes domum viderunt puerum cum Maria matre eius, et procidentes adoraverunt eum; et apertis thesauris suis, obtulerunt ei munera, aurum et tus et myrrham.
MATT|2|12|Et responso accepto in somnis, ne redirent ad Herodem, per aliam viam reversi sunt in regionem suam.
MATT|2|13|Qui cum recessissent, ecce angelus Domini apparet in somnis Ioseph dicens: " Surge et accipe puerum et matrem eius et fuge in Aegyptum et esto ibi, usque dum dicam tibi; futurum est enim ut Herodes quaerat puerum ad perdendum eum ".
MATT|2|14|Qui consurgens accepit puerum et matrem eius nocte et recessit in Aegyptum
MATT|2|15|et erat ibi usque ad obitum Herodis, ut adimpleretur, quod dictum est a Domino per prophetam dicentem: Ex Aegypto vocavi filium meum ".
MATT|2|16|Tunc Herodes videns quoniam illusus esset a Magis, iratus est valde et mittens occidit omnes pueros, qui erant in Bethlehem et in omnibus finibus eius, a bimatu et infra, secundum tempus, quod exquisierat a Magis.
MATT|2|17|Tunc adimpletum est, quod dictum est per Ieremiam prophetam dicentem:
MATT|2|18|" Vox in Rama audita est,ploratus et ululatus multus:Rachel plorans filios suos,et noluit consolari, quia non sunt ".
MATT|2|19|Defuncto autem Herode, ecce apparet angelus Domini in somnis Ioseph in Aegypto
MATT|2|20|dicens: " Surge et accipe puerum et matrem eius et vade in terram Israel; defuncti sunt enim, qui quaerebant animam pueri ".
MATT|2|21|Qui surgens accepit puerum et matrem eius et venit in terram Israel.
MATT|2|22|Audiens autem quia Archelaus regnaret in Iudaea pro Herode patre suo, timuit illuc ire; et admonitus in somnis, secessit in partes Galilaeae
MATT|2|23|et veniens habitavit in civitate, quae vocatur Nazareth, ut adimpleretur, quod dictum est per Prophetas: " Nazaraeus vocabitur ".
MATT|3|1|In diebus autem illis venit Ioannes Baptista praedicans in deserto Iudaeae
MATT|3|2|et dicens: " Paenitentiam agite; appropinquavit enim regnum caelorum ".
MATT|3|3|Hic est enim, qui dictus est per Isaiam prophetam dicentem: Vox clamantis in deserto:Parate viam Domini,rectas facite semitas eius!" ".
MATT|3|4|Ipse autem Ioannes habebat vestimentum de pilis cameli et zonam pelliceam circa lumbos suos; esca autem eius erat locustae et mel silvestre.
MATT|3|5|Tunc exibat ad eum Hierosolyma et omnis Iudaea et omnis regio circa Iordanem,
MATT|3|6|et baptizabantur in Iordane flumine ab eo, confitentes peccata sua.
MATT|3|7|Videns autem multos pharisaeorum et sadducaeorum venientes ad baptismum suum, dixit eis: " Progenies viperarum, quis demonstravit vobis fugere a futura ira?
MATT|3|8|Facite ergo fructum dignum paenitentiae
MATT|3|9|et ne velitis dicere intra vos: "Patrem habemus Abraham"; dico enim vobis quoniam potest Deus de lapidibus istis suscitare Abrahae filios.
MATT|3|10|Iam enim securis ad radicem arborum posita est; omnis ergo arbor, quae non facit fructum bonum, exciditur et in ignem mittitur.
MATT|3|11|Ego quidem vos baptizo in aqua in paenitentiam; qui autem post me venturus est, fortior me est, cuius non sum dignus calceamenta portare; ipse vos baptizabit in Spiritu Sancto et igni,
MATT|3|12|cuius ventilabrum in manu sua, et permundabit aream suam et congregabit triticum suum in horreum, paleas autem comburet igni inexstinguibili ".
MATT|3|13|Tunc venit Iesus a Galilaea in Iordanem ad Ioannem, ut baptizaretur ab eo.
MATT|3|14|Ioannes autem prohibebat eum dicens: " Ego a te debeo baptizari, et tu venis ad me? ".
MATT|3|15|Respondens autem Iesus dixit ei: " Sine modo, sic enim decet nos implere omnem iustitiam ". Tunc dimittit eum.
MATT|3|16|Baptizatus autem Iesus, confestim ascendit de aqua; et ecce aperti sunt ei caeli, et vidit Spiritum Dei descendentem sicut columbam et venientem super se.
MATT|3|17|Et ecce vox de caelis dicens: "Hic est Filius meus dilectus, in quomihi complacui ".
MATT|4|1|Tunc Iesus ductus est in de sertum a Spiritu, ut tentaretur a Diabolo.
MATT|4|2|Et cum ieiunasset quadraginta diebus et quadraginta noctibus, postea esuriit.
MATT|4|3|Et accedens tentator dixit ei: " Si Filius Dei es, dic, ut lapides isti panes fiant ".
MATT|4|4|Qui respondens dixit: Scriptum est:Non in pane solo vivet homo,sed in omni verbo, quod procedit de ore Dei" ".
MATT|4|5|Tunc assumit eum Diabolus in sanctam civitatem et statuit eum supra pinnaculum templi
MATT|4|6|et dicit ei: " Si Filius Dei es, mitte te deorsum. Scriptum est enim:Angelis suis mandabit de te,et in manibus tollent te,ne forte offendas ad lapidem pedem tuum" ".
MATT|4|7|Ait illi Iesus: " Rursum scriptum est: "Non tentabis Dominum Deum tuum".
MATT|4|8|Iterum assumit eum Diabolus in montem excelsum valde et ostendit ei omnia regna mundi et gloriam eorum
MATT|4|9|et dicit illi: " Haec tibi omnia dabo, si cadens adoraveris me".
MATT|4|10|Tunc dicit ei Iesus: Vade, Satanas! Scriptum est enim:Dominum Deum tuum adorabiset illi soli servies" ".
MATT|4|11|Tunc reliquit eum Diabolus, et ecce angeli accesserunt et ministrabant ei.
MATT|4|12|Cum autem audisset quod Ioannes traditus esset, secessit in Galilaeam.
MATT|4|13|Et relicta Nazareth, venit et habitavit in Capharnaum maritimam
MATT|4|14|in finibus Zabulon et Nephthali, ut impleretur, quod dictum est per Isaiam prophetam dicentem:
MATT|4|15|" Terra Zabulon et terra Nephthali,ad viam maris, trans Iordanem,Galilaea gentium;
MATT|4|16|populus, qui sedebat in tenebris,lucem vidit magnam,et sedentibus in regione et umbra mortislux orta est eis ".
MATT|4|17|Exinde coepit Iesus praedicare et dicere: " Paenitentiam agite; appropinquavit enim regnum caelorum ".
MATT|4|18|Ambulans autem iuxta mare Galilaeae, vidit duos fratres, Simonem, qui vocatur Petrus, et Andream fratrem eius, mittentes rete in mare; erant enim piscatores.
MATT|4|19|Et ait illis: " Venite post me, et faciam vos piscatores hominum ".
MATT|4|20|At illi continuo, relictis retibus, secuti sunt eum.
MATT|4|21|Et procedens inde vidit alios duos fratres, Iacobum Zebedaei et Ioannem fratrem eius, in navi cum Zebedaeo patre eorum reficientes retia sua; et vocavit eos.
MATT|4|22|Illi autem statim, relicta navi et patre suo, secuti sunt eum.
MATT|4|23|Et circumibat Iesus totam Galilaeam, docens in synagogis eorum et praedicans evangelium regni et sanans omnem languorem et omnem infirmitatem in populo.
MATT|4|24|Et abiit opinio eius in totam Syriam; et obtulerunt ei omnes male habentes, variis languoribus et tormentis comprehensos, et qui daemonia habebant, et lunaticos et paralyticos, et curavit eos.
MATT|4|25|Et secutae sunt eum turbae multae de Galilaea et Decapoli et Hierosolymis et Iudaea et de trans Iordanem.
MATT|5|1|Videns autem turbas, ascendit in montem; et cum sedisset, ac cesserunt ad eum discipuli eius;
MATT|5|2|et aperiens os suum docebat eos dicens:
MATT|5|3|" Beati pauperes spiritu, quoniam ipsorum est regnum caelorum.
MATT|5|4|Beati, qui lugent, quoniam ipsi consolabuntur.
MATT|5|5|Beati mites, quoniam ipsi possidebunt terram.
MATT|5|6|Beati, qui esuriunt et sitiunt iustitiam, quoniam ipsi saturabuntur.
MATT|5|7|Beati misericordes, quia ipsi misericordiam consequentur.
MATT|5|8|Beati mundo corde, quoniam ipsi Deum videbunt.
MATT|5|9|Beati pacifici, quoniam filii Dei vocabuntur.
MATT|5|10|Beati, qui persecutionem patiuntur propter iustitiam, quoniam ipsorum est regnum caelorum.
MATT|5|11|Beati estis cum maledixerint vobis et persecuti vos fuerint et dixerint omne malum adversum vos, mentientes, propter me.
MATT|5|12|Gaudete et exsultate, quoniam merces vestra copiosa est in caelis; sic enim persecuti sunt prophetas, qui fuerunt ante vos.
MATT|5|13|Vos estis sal terrae; quod si sal evanuerit, in quo salietur? Ad nihilum valet ultra, nisi ut mittatur foras et conculcetur ab hominibus.
MATT|5|14|Vos estis lux mundi. Non potest civitas abscondi supra montem posita;
MATT|5|15|neque accendunt lucernam et ponunt eam sub modio, sed super candelabrum, ut luceat omnibus, qui in domo sunt.
MATT|5|16|Sic luceat lux vestra coram hominibus, ut videant vestra bona opera et glorificent Patrem vestrum, qui in caelis est.
MATT|5|17|Nolite putare quoniam veni solvere Legem aut Prophetas; non veni solvere, sed adimplere.
MATT|5|18|Amen quippe dico vobis: Donec transeat caelum et terra, iota unum aut unus apex non praeteribit a Lege, donec omnia fiant.
MATT|5|19|Qui ergo solverit unum de mandatis istis minimis et docuerit sic homines, minimus vocabitur in regno caelorum; qui autem fecerit et docuerit, hic magnus vocabitur in regno caelorum.
MATT|5|20|Dico enim vobis: Nisi abundaverit iustitia vestra plus quam scribarum et pharisaeorum, non intrabitis in regnum caelorum.
MATT|5|21|Audistis quia dictum est antiquis: "Non occides; qui autem occiderit, reus erit iudicio".
MATT|5|22|Ego autem dico vobis: Omnis, qui irascitur fratri suo, reus erit iudicio; qui autem dixerit fratri suo: "Racha", reus erit concilio; qui autem dixerit: "Fatue", reus erit gehennae ignis.
MATT|5|23|Si ergo offeres munus tuum ad altare, et ibi recordatus fueris quia frater tuus habet aliquid adversum te,
MATT|5|24|relinque ibi munus tuum ante altare et vade, prius, reconciliare fratri tuo et tunc veniens offer munus tuum.
MATT|5|25|Esto consentiens adversario tuo cito, dum es in via cum eo, ne forte tradat te adversarius iudici, et iudex tradat te ministro, et in carcerem mittaris.
MATT|5|26|Amen dico tibi: Non exies inde, donec reddas novissimum quadrantem.
MATT|5|27|Audistis quia dictum est: "Non moechaberis".
MATT|5|28|Ego autem dico vobis: Omnis, qui viderit mulierem ad concupiscendum eam, iam moechatus est eam in corde suo.
MATT|5|29|Quod si oculus tuus dexter scandalizat te, erue eum et proice abs te; expedit enim tibi, ut pereat unum membrorum tuorum, quam totum corpus tuum mittatur in gehennam.
MATT|5|30|Et si dextera manus tua scandalizat te, abscide eam et proice abs te; expedit enim tibi, ut pereat unum membrorum tuorum, quam totum corpus tuum abeat in gehennam.
MATT|5|31|Dictum est autem: "Quicumque dimiserit uxorem suam, det illi libellum repudii".
MATT|5|32|Ego autem dico vobis: Omnis, qui dimiserit uxorem suam, excepta fornicationis causa, facit eam moechari; et, qui dimissam duxerit, adulterat.
MATT|5|33|Iterum audistis quia dictum est antiquis: "Non periurabis; reddes autem Domino iuramenta tua".
MATT|5|34|Ego autem dico vobis: Non iurare omnino, neque per caelum, quia thronus Dei est,
MATT|5|35|neque per terram, quia scabellum est pedum eius, neque per Hierosolymam, quia civitas est magni Regis;
MATT|5|36|neque per caput tuum iuraveris, quia non potes unum capillum album facere aut nigrum.
MATT|5|37|Sit autem sermo vester: "Est, est", "Non, non"; quod autem his abundantius est, a Malo est.
MATT|5|38|Audistis quia dictum est: "Oculum pro oculo et dentem pro dente".
MATT|5|39|Ego autem dico vobis: Non resistere malo; sed si quis te percusserit in dextera maxilla tua, praebe illi et alteram;
MATT|5|40|et ei, qui vult tecum iudicio contendere et tunicam tuam tollere, remitte ei et pallium;
MATT|5|41|et quicumque te angariaverit mille passus, vade cum illo duo.
MATT|5|42|Qui petit a te, da ei; et volenti mutuari a te, ne avertaris.
MATT|5|43|Audistis quia dictum est: "Diliges proximum tuum et odio habebis inimicum tuum".
MATT|5|44|Ego autem dico vobis: Diligite inimicos vestros et orate pro persequentibus vos,
MATT|5|45|ut sitis filii Patris vestri, qui in caelis est, quia solem suum oriri facit super malos et bonos et pluit super iustos et iniustos.
MATT|5|46|Si enim dilexeritis eos, qui vos diligunt, quam mercedem habetis? Nonne et publicani hoc faciunt?
MATT|5|47|Et si salutaveritis fratres vestros tantum, quid amplius facitis? Nonne et ethnici hoc faciunt?
MATT|5|48|Estote ergo vos perfecti, sicut Pater vester caelestis perfectus est.
MATT|6|1|Attendite, ne iustitiam vestram faciatis coram hominibus, ut vi deamini ab eis; alioquin mercedem non habetis apud Patrem vestrum, qui in caelis est.
MATT|6|2|Cum ergo facies eleemosynam, noli tuba canere ante te, sicut hypocritae faciunt in synagogis et in vicis, ut honorificentur ab hominibus. Amen dico vobis: Receperunt mercedem suam.
MATT|6|3|Te autem faciente eleemosynam, nesciat sinistra tua quid faciat dextera tua,
MATT|6|4|ut sit eleemosyna tua in abscondito, et Pater tuus, qui videt in abscondito, reddet tibi.
MATT|6|5|Et cum oratis, non eritis sicut hypocritae, qui amant in synagogis et in angulis platearum stantes orare, ut videantur ab hominibus. Amen dico vobis: Receperunt mercedem suam.
MATT|6|6|Tu autem cum orabis, intra in cubiculum tuum et, clauso ostio tuo, ora Patrem tuum, qui est in abscondito; et Pater tuus, qui videt in abscondito, reddet tibi.
MATT|6|7|Orantes autem nolite multum loqui sicut ethnici; putant enim quia in multiloquio suo exaudiantur.
MATT|6|8|Nolite ergo assimilari eis; scit enim Pater vester, quibus opus sit vobis, antequam petatis eum.
MATT|6|9|Sic ergo vos orabitis:Pater noster, qui es in caelis,sanctificetur nomen tuum,
MATT|6|10|adveniat regnum tuum,fiat voluntas tua,sicut in caelo, et in terra.
MATT|6|11|Panem nostrum supersubstantialem da nobis hodie;
MATT|6|12|et dimitte nobis debita nostra,sicut et nos dimittimus debitoribus nostris;
MATT|6|13|et ne inducas nos in tentationem,sed libera nos a Malo.
MATT|6|14|Si enim dimiseritis hominibus peccata eorum, dimittet et vobis Pater vester caelestis;
MATT|6|15|si autem non dimiseritis hominibus, nec Pater vester dimittet peccata vestra.
MATT|6|16|Cum autem ieiunatis, nolite fieri sicut hypocritae tristes; demoliuntur enim facies suas, ut pareant hominibus ieiunantes. Amen dico vobis: Receperunt mercedem suam.
MATT|6|17|Tu autem cum ieiunas, unge caput tuum et faciem tuam lava,
MATT|6|18|ne videaris hominibus ieiunans sed Patri tuo, qui est in abscondito; et Pater tuus, qui videt in abscondito, reddet tibi.
MATT|6|19|Nolite thesaurizare vobis thesauros in terra, ubi aerugo et tinea demolitur, et ubi fures effodiunt et furantur;
MATT|6|20|thesaurizate autem vobis thesauros in caelo, ubi neque aerugo neque tinea demolitur, et ubi fures non effodiunt nec furantur;
MATT|6|21|ubi enim est thesaurus tuus, ibi erit et cor tuum.
MATT|6|22|Lucerna corporis est oculus. Si ergo fuerit oculus tuus simplex, totum corpus tuum lucidum erit;
MATT|6|23|si autem oculus tuus nequam fuerit, totum corpus tuum tenebrosum erit. Si ergo lumen, quod in te est, tene brae sunt, tenebrae quantae erunt!
MATT|6|24|Nemo potest duobus dominis servire: aut enim unum odio habebit et alterum diliget, aut unum sustinebit et alterum contemnet; non potestis Deo servire et mammonae.
MATT|6|25|Ideo dico vobis: Ne solliciti sitis animae vestrae quid manducetis, neque corpori vestro quid induamini. Nonne anima plus est quam esca, et corpus quam vestimentum?
MATT|6|26|Respicite volatilia caeli, quoniam non serunt neque metunt neque congregant in horrea, et Pater vester caelestis pascit illa. Nonne vos magis pluris estis illis?
MATT|6|27|Quis autem vestrum cogitans potest adicere ad aetatem suam cubitum unum?
MATT|6|28|Et de vestimento quid solliciti estis? Considerate lilia agri quomodo crescunt: non laborant neque nent.
MATT|6|29|Dico autem vobis quoniam nec Salomon in omni gloria sua coopertus est sicut unum ex istis.
MATT|6|30|Si autem fenum agri, quod hodie est et cras in clibanum mittitur, Deus sic vestit, quanto magis vos, modicae fidei?
MATT|6|31|Nolite ergo solliciti esse dicentes: "Quid manducabimus?", aut: "Quid bibemus?", aut: "Quo operiemur?".
MATT|6|32|Haec enim omnia gentes inquirunt; scit enim Pater vester caelestis quia his omnibus indigetis.
MATT|6|33|Quaerite autem primum regnum Dei et iustitiam eius, et haec omnia adicientur vobis.
MATT|6|34|Nolite ergo esse solliciti in crastinum; crastinus enim dies sollicitus erit sibi ipse. Sufficit diei malitia sua.
MATT|7|1|Nolite iudicare, ut non iudice mini;
MATT|7|2|in quo enim iudicio iudi caveritis, iudicabimini, et in qua mensura mensi fueritis, metietur vobis.
MATT|7|3|Quid autem vides festucam in oculo fratris tui, et trabem in oculo tuo non vides?
MATT|7|4|Aut quomodo dices fratri tuo: "Sine, eiciam festucam de oculo tuo", et ecce trabes est in oculo tuo?
MATT|7|5|Hypocrita, eice primum trabem de oculo tuo, et tunc videbis eicere festucam de oculo fratris tui.
MATT|7|6|Nolite dare sanctum canibus neque mittatis margaritas vestras ante porcos, ne forte conculcent eas pedibus suis et conversi dirumpant vos.
MATT|7|7|Petite, et dabitur vobis; quaerite et invenietis; pulsate, et aperietur vobis.
MATT|7|8|Omnis enim qui petit, accipit; et, qui quaerit, invenit; et pulsanti aperietur.
MATT|7|9|Aut quis est ex vobis homo, quem si petierit filius suus panem, numquid lapidem porriget ei?
MATT|7|10|Aut si piscem petierit, numquid serpentem porriget ei?
MATT|7|11|Si ergo vos, cum sitis mali, nostis dona bona dare filiis vestris, quanto magis Pater vester, qui in caelis est, dabit bona petentibus se.
MATT|7|12|Omnia ergo, quaecumque vultis ut faciant vobis homines, ita et vos facite eis; haec est enim Lex et Prophetae.
MATT|7|13|Intrate per angustam portam, quia lata porta et spatiosa via, quae ducit ad perditionem, et multi sunt, qui intrant per eam;
MATT|7|14|quam angusta porta et arta via, quae ducit ad vitam, et pauci sunt, qui inveniunt eam!
MATT|7|15|Attendite a falsis prophetis, qui veniunt ad vos in vestimentis ovium, intrinsecus autem sunt lupi rapaces.
MATT|7|16|A fructibus eorum cognoscetis eos; numquid colligunt de spinis uvas aut de tribulis ficus?
MATT|7|17|Sic omnis arbor bona fructus bonos facit, mala autem arbor fructus malos facit;
MATT|7|18|non potest arbor bona fructus malos facere, neque arbor mala fructus bonos facere.
MATT|7|19|Omnis arbor, quae non facit fructum bonum, exciditur et in ignem mittitur.
MATT|7|20|Igitur ex fructibus eorum cognoscetis eos.
MATT|7|21|Non omnis, qui dicit mihi: "Domine, Domine", intrabit in regnum caelorum, sed qui facit voluntatem Patris mei, qui in caelis est.
MATT|7|22|Multi dicent mihi in illa die: "Domine, Domine, nonne in tuo nomine prophetavimus, et in tuo nomine daemonia eiecimus, et in tuo nomine virtutes multas fecimus?".
MATT|7|23|Et tunc confitebor illis: Numquam novi vos; discedite a me, qui operamini iniquitatem.
MATT|7|24|Omnis ergo, qui audit verba mea haec et facit ea, assimilabitur viro sapienti, qui aedificavit domum suam supra petram.
MATT|7|25|Et descendit pluvia, et venerunt flumina, et flaverunt venti et irruerunt in domum illam, et non cecidit; fundata enim erat supra petram.
MATT|7|26|Et omnis, qui audit verba mea haec et non facit ea, similis erit viro stulto, qui aedificavit domum suam supra arenam.
MATT|7|27|Et descendit pluvia, et venerunt flumina, et flaverunt venti et irruerunt in domum illam, et cecidit, et fuit ruina eius magna ".
MATT|7|28|Et factum est, cum consummasset Iesus verba haec, admirabantur turbae super doctrinam eius;
MATT|7|29|erat enim docens eos sicut potestatem habens, et non sicut scribae eorum.
MATT|8|1|Cum autem descendisset de monte, secutae sunt eum turbae multae.
MATT|8|2|Et ecce leprosus veniens adorabat eum dicens: " Domine, si vis, potes me mundare ".
MATT|8|3|Et extendens manum, tetigit eum dicens: " Volo, mundare! "; et confestim mundata est lepra eius.
MATT|8|4|Et ait illi Iesus: " Vide, nemini dixeris; sed vade, ostende te sacerdoti et offer munus, quod praecepit Moyses, in testimonium illis ".
MATT|8|5|Cum autem introisset Capharnaum, accessit ad eum centurio rogans eum
MATT|8|6|et dicens: " Domine, puer meus iacet in domo paralyticus et male torquetur ".
MATT|8|7|Et ait illi: " Ego veniam et curabo eum ".
MATT|8|8|Et respondens centurio ait: " Domine, non sum dignus, ut intres sub tectum meum, sed tantum dic verbo, et sanabitur puer meus.
MATT|8|9|Nam et ego homo sum sub potestate, habens sub me milites, et dico huic: Vade", et vadit; et alii: "Veni", et venit; et servo meo: "Fac hoc", et facit".
MATT|8|10|Audiens autem Iesus, miratus est et sequentibus se dixit: "Amen dico vobis: Apud nullum inveni tantam fidem in Israel!
MATT|8|11|Dico autem vobis quod multi ab oriente et occidente venient et recumbent cum Abraham et Isaac et Iacob in regno caelorum;
MATT|8|12|filii autem regni eicientur in tenebras exteriores: ibi erit fletus et stridor dentium ".
MATT|8|13|Et dixit Iesus centurioni: " Vade; sicut credidisti, fiat tibi ". Et sanatus est puer in hora illa.
MATT|8|14|Et cum venisset Iesus in domum Petri, vidit socrum eius iacentem et febricitantem;
MATT|8|15|et tetigit manum eius, et dimisit eam febris; et surrexit et ministrabat ei.
MATT|8|16|Vespere autem facto, obtulerunt ei multos daemonia habentes; et eiciebat spiritus verbo et omnes male habentes curavit,
MATT|8|17|ut adimpleretur, quod dictum est per Isaiam prophetam dicentem: Ipse infirmitates nostras accepitet aegrotationes portavit ".
MATT|8|18|Videns autem Iesus turbas multas circum se, iussit ire trans fretum.
MATT|8|19|Et accedens unus scriba ait illi: " Magister, sequar te, quocumque ieris ".
MATT|8|20|Et dicit ei Iesus: " Vulpes foveas habent, et volucres caeli tabernacula, Filius autem hominis non habet, ubi caput reclinet ".
MATT|8|21|Alius autem de discipulis eius ait illi: "Domine, permitte me primum ire et sepelire patrem meum ".
MATT|8|22|Iesus autem ait illi: " Sequere me et dimitte mortuos sepelire mortuos suos ".
MATT|8|23|Et ascendente eo in naviculam, secuti sunt eum discipuli eius.
MATT|8|24|Et ecce motus magnus factus est in mari, ita ut navicula operiretur fluctibus; ipse vero dormiebat.
MATT|8|25|Et accesserunt et suscitaverunt eum dicentes: " Domine, salva nos, perimus! ".
MATT|8|26|Et dicit eis: " Quid timidi estis, modicae fidei? ". Tunc surgens increpavit ventis et mari, et facta est tranquillitas magna.
MATT|8|27|Porro homines mirati sunt dicentes: " Qualis est hic, quia et venti et mare oboediunt ei? ".
MATT|8|28|Et cum venisset trans fretum in regionem Gadarenorum, occurrerunt ei duo habentes daemonia, de monumentis exeuntes, saevi nimis, ita ut nemo posset transire per viam illam.
MATT|8|29|Et ecce clamaverunt dicentes: " Quid nobis et tibi, Fili Dei? Venisti huc ante tempus torquere nos? ".
MATT|8|30|Erat autem longe ab illis grex porcorum multorum pascens.
MATT|8|31|Daemones autem rogabant eum dicentes: " Si eicis nos, mitte nos in gregem porcorum ".
MATT|8|32|Et ait illis: " Ite ". Et illi exeuntes abierunt in porcos; et ecce impetu abiit totus grex per praeceps in mare, et mortui sunt in aquis.
MATT|8|33|Pastores autem fugerunt et venientes in civitatem nuntiaverunt omnia et de his, qui daemonia habuerant.
MATT|8|34|Et ecce tota civitas exiit obviam Iesu, et viso eo rogabant, ut transiret a finibus eorum.
MATT|9|1|Et ascendens in naviculam transfretavit et venit in civita tem suam.
MATT|9|2|Et ecce offerebant ei paralyticum iacentem in lecto. Et videns Iesus fidem illorum, dixit paralytico: " Confide, fili; remittuntur peccata tua.
MATT|9|3|Et ecce quidam de scribis dixerunt intra se: " Hic blasphemat ".
MATT|9|4|Et cum vidisset Iesus cogitationes eorum, dixit: " Ut quid cogitatis mala in cordibus vestris?
MATT|9|5|Quid enim est facilius, dicere: "Dimittuntur peccata tua", aut dicere: Surge et ambula"?
MATT|9|6|Ut sciatis autem quoniam Filius hominis habet potestatem in terra dimittendi peccata - tunc ait paralytico -: Surge, tolle lectum tuum et vade in domum tuam ".
MATT|9|7|Et surrexit et abiit in domum suam.
MATT|9|8|Videntes autem turbae timuerunt et glorificaverunt Deum, qui dedit potestatem talem hominibus.
MATT|9|9|Et cum transiret inde Iesus, vidit hominem sedentem in teloneo, Matthaeum nomine, et ait illi: "Sequere me". Et surgens secutus est eum.
MATT|9|10|Et factum est, discumbente eo in domo, ecce multi publicani et peccatores venientes simul discumbebant cum Iesu et discipulis eius.
MATT|9|11|Et videntes pharisaei dicebant discipulis eius: " Quare cum publicanis et peccatoribus manducat magister vester? ".
MATT|9|12|At ille audiens ait: " Non est opus valentibus medico sed male habentibus.
MATT|9|13|Euntes autem discite quid est: "Misericordiam volo et non sacrificium". Non enim veni vocare iustos sed peccatores ".
MATT|9|14|Tunc accedunt ad eum discipuli Ioannis dicentes: " Quare nos et pharisaei ieiunamus frequenter, discipuli autem tui non ieiunant? ".
MATT|9|15|Et ait illis Iesus: " Numquid possunt convivae nuptiarum lugere, quamdiu cum illis est sponsus? Venient autem dies, cum auferetur ab eis sponsus, et tunc ieiunabunt.
MATT|9|16|Nemo autem immittit commissuram panni rudis in vestimentum vetus; tollit enim supplementum eius a vestimento, et peior scissura fit.
MATT|9|17|Neque mittunt vinum novum in utres veteres, alioquin rumpuntur utres, et vinum effunditur, et utres pereunt; sed vinum novum in utres novos mittunt, et ambo conservantur ".
MATT|9|18|Haec illo loquente ad eos, ecce princeps unus accessit et adorabat eum dicens: " Filia mea modo defuncta est; sed veni, impone manum tuam super eam, et vivet ".
MATT|9|19|Et surgens Iesus sequebatur eum et discipuli eius.
MATT|9|20|Et ecce mulier, quae sanguinis fluxum patiebatur duodecim annis, accessit retro et tetigit fimbriam vestimenti eius.
MATT|9|21|Dicebat enim intra se: " Si tetigero tantum vestimentum eius, salva ero.
MATT|9|22|At Iesus conversus et videns eam dixit: " Confide, filia; fides tua te salvam fecit ". Et salva facta est mulier ex illa hora.
MATT|9|23|Et cum venisset Iesus in domum principis et vidisset tibicines et turbam tumultuantem,
MATT|9|24|dicebat: " Recedite; non est enim mortua puella, sed dormit ". Et deridebant eum.
MATT|9|25|At cum eiecta esset turba, intravit et tenuit manum eius, et surrexit puella.
MATT|9|26|Et exiit fama haec in universam terram illam.
MATT|9|27|Et transeunte inde Iesu, secuti sunt eum duo caeci clamantes et dicentes: " Miserere nostri, fili David! ".
MATT|9|28|Cum autem venisset domum, accesserunt ad eum caeci, et dicit eis Iesus: Creditis quia possum hoc facere? ". Dicunt ei: "Utique, Domine".
MATT|9|29|Tunc tetigit oculos eorum dicens: "Secundum fidem vestram fiat vobis".
MATT|9|30|Et aperti sunt oculi illorum. Et comminatus est illis Iesus dicens: " Videte, ne quis sciat ".
MATT|9|31|Illi autem exeuntes diffamaverunt eum in universa terra illa.
MATT|9|32|Egressis autem illis, ecce obtulerunt ei hominem mutum, daemonium habentem.
MATT|9|33|Et eiecto daemone, locutus est mutus. Et miratae sunt turbae dicentes: Numquam apparuit sic in Israel! ".
MATT|9|34|Pharisaei autem dicebant: " In principe daemoniorum eicit daemones ".
MATT|9|35|Et circumibat Iesus civitates omnes et castella, docens in synagogis eorum et praedicans evangelium regni et curans omnem languorem et omnem infirmitatem.
MATT|9|36|Videns autem turbas, misertus est eis, quia erant vexati et iacentes sicut oves non habentes pastorem.
MATT|9|37|Tunc dicit discipulis suis: " Messis quidem multa, operarii autem pauci;
MATT|9|38|rogate ergo Dominum messis, ut mittat operarios in messem suam ".
MATT|10|1|Et convocatis Duodecim di scipulis suis, dedit illis pote statem spirituum immundorum, ut eicerent eos et curarent omnem languorem et omnem infirmitatem.
MATT|10|2|Duodecim autem apostolorum nomina sunt haec: primus Simon, qui dicitur Petrus, et Andreas frater eius, et Iacobus Zebedaei et Ioannes frater eius,
MATT|10|3|Philippus et Bartholomaeus, Thomas et Matthaeus publicanus, Iacobus Alphaei et Thaddaeus,
MATT|10|4|Simon Chananaeus et Iudas Iscariotes, qui et tradidit eum.
MATT|10|5|Hos Duodecim misit Iesus praecipiens eis et dicens: " In viam gentium ne abieritis et in civitates Samaritanorum ne intraveritis;
MATT|10|6|sed potius ite ad oves, quae perierunt domus Israel.
MATT|10|7|Euntes autem praedicate dicentes: "Appropinquavit regnum caelorum".
MATT|10|8|Infirmos curate, mortuos suscitate, leprosos mundate, daemones eicite; gratis accepistis, gratis date.
MATT|10|9|Nolite possidere aurum neque argentum neque pecuniam in zonis vestris,
MATT|10|10|non peram in via neque duas tunicas neque calceamenta neque virgam; dignus enim est operarius cibo suo.
MATT|10|11|In quamcumque civitatem aut castellum intraveritis, interrogate quis in ea dignus sit; et ibi manete donec exeatis.
MATT|10|12|Intrantes autem in domum, salutate eam;
MATT|10|13|et si quidem fuerit domus digna, veniat pax vestra super eam; si autem non fuerit digna, pax vestra ad vos revertatur.
MATT|10|14|Et quicumque non receperit vos neque audierit sermones vestros, exeuntes foras de domo vel de civitate illa, excutite pulverem de pedibus vestris.
MATT|10|15|Amen dico vobis: Tolerabilius erit terrae Sodomorum et Gomorraeorum in die iudicii quam illi civitati.
MATT|10|16|Ecce ego mitto vos sicut oves in medio luporum; estote ergo prudentes sicut serpentes et simplices sicut columbae.
MATT|10|17|Cavete autem ab hominibus; tradent enim vos in conciliis, et in synagogis suis flagellabunt vos;
MATT|10|18|et ad praesides et ad reges ducemini propter me in testimonium illis et gentibus.
MATT|10|19|Cum autem tradent vos, nolite cogitare quomodo aut quid loquamini; dabitur enim vobis in illa hora quid loquamini.
MATT|10|20|Non enim vos estis, qui loquimini, sed Spiritus Patris vestri, qui loquitur in vobis.
MATT|10|21|Tradet autem frater fratrem in mortem, et pater filium; et insurgent filii in parentes et morte eos afficient.
MATT|10|22|Et eritis odio omnibus propter nomen meum; qui autem perseveraverit in finem, hic salvus erit.
MATT|10|23|Cum autem persequentur vos in civitate ista, fugite in aliam; amen enim dico vobis: Non consummabitis civitates Israel, donec veniat Filius hominis.
MATT|10|24|Non est discipulus super magistrum nec servus super dominum suum.
MATT|10|25|Sufficit discipulo, ut sit sicut magister eius, et servus sicut dominus eius. Si patrem familias Beelzebul vocaverunt, quanto magis domesticos eius!
MATT|10|26|Ne ergo timueritis eos. Nihil enim est opertum, quod non revelabitur, et occultum, quod non scietur.
MATT|10|27|Quod dico vobis in tenebris, dicite in lumine; et, quod in aure auditis, praedicate super tecta.
MATT|10|28|Et nolite timere eos, qui occidunt corpus, animam autem non possunt occidere; sed potius eum timete, qui potest et animam et corpus perdere in gehenna.
MATT|10|29|Nonne duo passeres asse veneunt? Et unus ex illis non cadet super terram sine Patre vestro.
MATT|10|30|Vestri autem et capilli capitis omnes numerati sunt.
MATT|10|31|Nolite ergo timere; multis passeribus meliores estis vos.
MATT|10|32|Omnis ergo qui confitebitur me coram hominibus, confitebor et ego eum coram Patre meo, qui est in caelis;
MATT|10|33|qui autem negaverit me coram hominibus, negabo et ego eum coram Patre meo, qui est in caelis.
MATT|10|34|Nolite arbitrari quia venerim mittere pacem in terram; non veni pacem mittere sed gladium.
MATT|10|35|Veni enim separarehominem adversus patrem suumet filiam adversus matrem suamet nurum adversus socrum suam:
MATT|10|36|et inimici hominis domestici eius.
MATT|10|37|Qui amat patrem aut matrem plus quam me, non est me dignus; et, qui amat filium aut filiam super me, non est me dignus;
MATT|10|38|et, qui non accipit crucem suam et sequitur me, non est me dignus.
MATT|10|39|Qui invenerit animam suam, perdet illam; et, qui perdiderit animam suam propter me, inveniet eam.
MATT|10|40|Qui recipit vos, me recipit; et, qui me recipit, recipit eum, qui me misit.
MATT|10|41|Qui recipit prophetam in nomine prophetae, mercedem prophetae accipiet; et, qui recipit iustum in nomine iusti, mercedem iusti accipiet.
MATT|10|42|Et, quicumque potum dederit uni ex minimis istis calicem aquae frigidae tantum in nomine discipuli, amen dico vobis: Non perdet mercedem suam ".
MATT|11|1|Et factum est, cum consum masset Iesus praecipiens Duodecim discipulis suis, transiit inde, ut doceret et praedicaret in civitatibus eorum.
MATT|11|2|Ioannes autem, cum audisset in vinculis opera Christi, mittens per discipulos suos
MATT|11|3|ait illi: " Tu es qui venturus es, an alium exspectamus? ".
MATT|11|4|Et respondens Iesus ait illis: " Euntes renuntiate Ioanni, quae auditis et videtis:
MATT|11|5|caeci vident et claudi ambulant, leprosi mundantur et surdi audiunt et mortui resurgunt et pauperes evangelizantur;
MATT|11|6|et beatus est, qui non fuerit scandalizatus in me ".
MATT|11|7|Illis autem abeuntibus, coepit Iesus dicere ad turbas de Ioanne: " Quid existis in desertum videre? Arundinem vento agitatam?
MATT|11|8|Sed quid existis videre? Hominem mollibus vestitum? Ecce, qui mollibus vestiuntur, in domibus regum sunt.
MATT|11|9|Sed quid existis videre? Prophetam? Etiam, dico vobis, et plus quam prophetam.
MATT|11|10|Hic est, de quo scriptum est:Ecce ego mitto angelum meum ante faciem tuam,qui praeparabit viam tuam ante te".
MATT|11|11|Amen dico vobis: Non surrexit inter natos mulierum maior Ioanne Baptista; qui autem minor est in regno caelorum, maior est illo.
MATT|11|12|A diebus autem Ioannis Baptistae usque nunc regnum caelorum vim patitur, et violenti rapiunt illud.
MATT|11|13|Omnes enim Prophetae et Lex usque ad Ioannem prophetaverunt;
MATT|11|14|et si vultis recipere, ipse est Elias, qui venturus est.
MATT|11|15|Qui habet aures, audiat.
MATT|11|16|Cui autem similem aestimabo generationem istam? Similis est pueris sedentibus in foro, qui clamantes coaequalibus
MATT|11|17|dicunt:Cecinimus vobis, et non saltastis;lamentavimus, et non planxistis".
MATT|11|18|Venit enim Ioannes neque manducans neque bibens, et dicunt: "Daemonium habet!";
MATT|11|19|venit Filius hominis manducans et bibens, et dicunt: "Ecce homo vorax et potator vini, publicanorum amicus et peccatorum!". Et iustificata est sapientia ab operibus suis ".
MATT|11|20|Tunc coepit exprobrare civitatibus, in quibus factae sunt plurimae virtutes eius, quia non egissent paenitentiam:
MATT|11|21|" Vae tibi, Chorazin! Vae tibi, Bethsaida! Quia si in Tyro et Sidone factae essent virtutes, quae factae sunt in vobis, olim in cilicio et cinere paenitentiam egissent.
MATT|11|22|Verumtamen dico vobis: Tyro et Sidoni remissius erit in die iudicii quam vobis.
MATT|11|23|Et tu, Capharnaum, numquid usque in caelum exaltaberis? Usque in infernum descendes! Quia si in Sodomis factae fuissent virtutes, quae factae sunt in te, mansissent usque in hunc diem.
MATT|11|24|Verumtamen dico vobis: Terrae Sodomorum remissius erit in die iudicii quam tibi ".
MATT|11|25|In illo tempore respondens Iesus dixit: " Confiteor tibi, Pater, Domine caeli et terrae, quia abscondisti haec a sapientibus et prudentibus et revelasti ea parvulis.
MATT|11|26|Ita, Pater, quoniam sic fuit placitum ante te.
MATT|11|27|Omnia mihi tradita sunt a Patre meo; et nemo novit Filium nisi Pater, neque Patrem quis novit nisi Filius et cui voluerit Filius revelare.
MATT|11|28|Venite ad me, omnes, qui laboratis et onerati estis, et ego reficiam vos.
MATT|11|29|Tollite iugum meum super vos et discite a me, quia mitis sum et humilis corde, et invenietis requiem animabus vestris.
MATT|11|30|Iugum enim meum suave, et onus meum leve est ".
MATT|12|1|In illo tempore abiit Iesus sabbatis per sata; discipuli autem eius esurierunt et coeperunt vellere spicas et manducare.
MATT|12|2|Pharisaei autem videntes dixerunt ei: " Ecce discipuli tui faciunt, quod non licet facere sabbato ".
MATT|12|3|At ille dixit eis: " Non legistis quid fecerit David, quando esuriit, et qui cum eo erant?
MATT|12|4|Quomodo intravit in domum Dei et panes propositionis comedit, quod non licebat ei edere neque his, qui cum eo erant, nisi solis sacerdotibus?
MATT|12|5|Aut non legistis in Lege quia sabbatis sacerdotes in templo sabbatum violant et sine crimine sunt?
MATT|12|6|Dico autem vobis quia templo maior est hic.
MATT|12|7|Si autem sciretis quid est: "Misericordiam volo et non sacrificium", numquam condemnassetis innocentes.
MATT|12|8|Dominus est enim Filius hominis sabbati ".
MATT|12|9|Et cum inde transisset, venit in synagogam eorum;
MATT|12|10|et ecce homo manum habens aridam. Et interrogabant eum dicentes: " Licet sabbatis curare? ", ut accusarent eum.
MATT|12|11|Ipse autem dixit illis: " Quis erit ex vobis homo, qui habeat ovem unam et, si ceciderit haec sabbatis in foveam, nonne tenebit et levabit eam?
MATT|12|12|Quanto igitur melior est homo ove! Itaque licet sabbatis bene facere ".
MATT|12|13|Tunc ait homini: " Extende manum tuam ". Et extendit, et restituta est sana sicut altera.
MATT|12|14|Exeuntes autem pharisaei consilium faciebant adversus eum, quomodo eum perderent.
MATT|12|15|Iesus autem sciens secessit inde. Et secuti sunt eum multi, et curavit eos omnes
MATT|12|16|et comminatus est eis, ne manifestum eum facerent,
MATT|12|17|ut adimpleretur, quod dictum est per Isaiam prophetam dicentem:
MATT|12|18|" Ecce puer meus, quem elegi,dilectus meus, in quo bene placuit animae meae;ponam Spiritum meum super eum,et iudicium gentibus nuntiabit.
MATT|12|19|Non contendet neque clamabit,neque audiet aliquis in plateis vocem eius.
MATT|12|20|Arundinem quassatam non confringetet linum fumigans non exstinguet,donec eiciat ad victoriam iudicium;
MATT|12|21|et in nomine eius gentes sperabunt ".
MATT|12|22|Tunc oblatus est ei daemonium habens, caecus et mutus, et curavit eum, ita ut mutus loqueretur et videret.
MATT|12|23|Et stupebant omnes turbae et dicebant: " Numquid hic est filius David?.
MATT|12|24|Pharisaei autem audientes dixerunt: " Hic non eicit daemones nisi in Beelzebul, principe daemonum ".
MATT|12|25|Sciens autem cogitationes eorum dixit eis: " Omne regnum divisum contra se desolatur, et omnis civitas vel domus divisa contra se non stabit.
MATT|12|26|Et si Satanas Satanam eicit, adversus se divisus est; quomodo ergo stabit regnum eius?
MATT|12|27|Et si ego in Beelzebul eicio daemones, filii vestri in quo eiciunt? Ideo ipsi iudices erunt vestri.
MATT|12|28|Si autem in Spiritu Dei ego eicio daemones, igitur pervenit in vos regnum Dei.
MATT|12|29|Aut quomodo potest quisquam intrare in domum fortis et vasa eius diripere, nisi prius alligaverit fortem? Et tunc domum illius diripiet.
MATT|12|30|Qui non est mecum, contra me est; et, qui non congregat mecum, spargit.
MATT|12|31|Ideo dico vobis: Omne peccatum et blasphemia remittetur hominibus, Spiritus autem blasphemia non remittetur.
MATT|12|32|Et quicumque dixerit verbum contra Filium hominis, remittetur ei; qui autem dixerit contra Spiritum Sanctum, non remittetur ei neque in hoc saeculo neque in futuro.
MATT|12|33|Aut facite arborem bonam et fructum eius bonum, aut facite arborem malam et fructum eius malum: si quidem ex fructu arbor agnoscitur.
MATT|12|34|Progenies viperarum, quomodo potestis bona loqui, cum sitis mali? Ex abundantia enim cordis os loquitur.
MATT|12|35|Bonus homo de bono thesauro profert bona, et malus homo de malo thesauro profert mala.
MATT|12|36|Dico autem vobis: Omne verbum otiosum, quod locuti fuerint homines, reddent rationem de eo in die iudicii:
MATT|12|37|ex verbis enim tuis iustificaberis, et ex verbis tuis condemnaberis ".
MATT|12|38|Tunc responderunt ei quidam de scribis et pharisaeis dicentes: " Magister, volumus a te signum videre ".
MATT|12|39|Qui respondens ait illis: " Generatio mala et adultera signum requirit; et signum non dabitur ei, nisi signum Ionae prophetae.
MATT|12|40|Sicut enim fuit Ionas in ventre ceti tribus diebus et tribus noctibus, sic erit Filius hominis in corde terrae tribus diebus et tribus noctibus.
MATT|12|41|Viri Ninevitae surgent in iudicio cum generatione ista et condemnabunt eam, quia paenitentiam egerunt in praedicatione Ionae; et ecce plus quam Iona hic!
MATT|12|42|Regina austri surget in iudicio cum generatione ista et condemnabit eam, quia venit a finibus terrae audire sapientiam Salomonis; et ecce plus quam Salomon hic!
MATT|12|43|Cum autem immundus spiritus exierit ab homine, ambulat per loca arida quaerens requiem et non invenit.
MATT|12|44|Tunc dicit: "Revertar in domum meam unde exivi"; et veniens invenit vacantem, scopis mundatam et ornatam.
MATT|12|45|Tunc vadit et assumit secum septem alios spiritus nequiores se, et intrantes habitant ibi; et fiunt novissima hominis illius peiora prioribus. Sic erit et generationi huic pessimae ".
MATT|12|46|Adhuc eo loquente ad turbas, ecce mater et fratres eius stabant foris quaerentes loqui ei.
MATT|12|47|Dixit autem ei quidam: " Ecce mater tua et fratres tui foris stant quaerentes loqui tecum ".
MATT|12|48|At ille respondens dicenti sibi ait: " Quae est mater mea, et qui sunt fratres mei? ".
MATT|12|49|Et extendens manum suam in discipulos suos dixit: " Ecce mater mea et fratres mei.
MATT|12|50|Quicumque enim fecerit voluntatem Patris mei, qui in caelis est, ipse meus frater et soror et mater est ".
MATT|13|1|In illo die exiens Iesus de domo sedebat secus mare;
MATT|13|2|et congregatae sunt ad eum turbae multae, ita ut in naviculam ascendens sederet, et omnis turba stabat in litore.
MATT|13|3|Et locutus est eis multa in parabolis dicens: " Ecce exiit, qui seminat, seminare.
MATT|13|4|Et dum seminat, quaedam ceciderunt secus viam, et venerunt volucres et comederunt ea.
MATT|13|5|Alia autem ceciderunt in petrosa, ubi non habebant terram multam, et continuo exorta sunt, quia non habebant altitudinem terrae;
MATT|13|6|sole autem orto, aestuaverunt et, quia non habebant radicem, aruerunt.
MATT|13|7|Alia autem ceciderunt in spinas, et creverunt spinae et suffocaverunt ea.
MATT|13|8|Alia vero ceciderunt in terram bonam et dabant fructum: aliud centesimum, aliud sexagesimum, aliud tricesimum.
MATT|13|9|Qui habet aures, audiat ".
MATT|13|10|Et accedentes discipuli dixerunt ei: " Quare in parabolis loqueris eis?.
MATT|13|11|Qui respondens ait illis: " Quia vobis datum est nosse mysteria regni caelorum, illis autem non est datum.
MATT|13|12|Qui enim habet, dabitur ei, et abundabit; qui autem non habet, et quod habet, auferetur ab eo.
MATT|13|13|Ideo in parabolis loquor eis, quia videntes non vident et audientes non audiunt neque intellegunt;
MATT|13|14|et adimpletur eis prophetia Isaiae dicens:Auditu audietis et non intellegetiset videntes videbitis et non videbitis.
MATT|13|15|Incrassatum est enim cor populi huius,et auribus graviter audieruntet oculos suos clauserunt,ne quando oculis videantet auribus audiantet corde intellegant et convertantur,et sanem eos".
MATT|13|16|Vestri autem beati oculi, quia vident, et aures vestrae, quia audiunt.
MATT|13|17|Amen quippe dico vobis: Multi prophetae et iusti cupierunt videre, quae videtis, et non viderunt, et audire, quae auditis, et non audierunt!
MATT|13|18|Vos ergo audite parabolam seminantis.
MATT|13|19|Omnis, qui audit verbum regni et non intellegit, venit Malus et rapit, quod seminatum est in corde eius; hic est, qui secus viam seminatus est.
MATT|13|20|Qui autem supra petrosa seminatus est, hic est, qui verbum audit et continuo cum gaudio accipit illud,
MATT|13|21|non habet autem in se radicem, sed est temporalis; facta autem tribulatione vel persecutione propter verbum, continuo scandalizatur.
MATT|13|22|Qui autem est seminatus in spinis, hic est, qui verbum audit, et sollicitudo saeculi et fallacia divitiarum suffocat verbum, et sine fructu efficitur.
MATT|13|23|Qui vero in terra bona seminatus est, hic est, qui audit verbum et intellegit et fructum affert et facit aliud quidem centum, aliud autem sexaginta, porro aliud triginta ".
MATT|13|24|Aliam parabolam proposuit illis dicens: " Simile factum est regnum caelorum homini, qui seminavit bonum semen in agro suo.
MATT|13|25|Cum autem dormirent homines, venit inimicus eius et superseminavit zizania in medio tritici et abiit.
MATT|13|26|Cum autem crevisset herba et fructum fecisset, tunc apparuerunt et zizania.
MATT|13|27|Accedentes autem servi patris familias dixerunt ei: "Domine, nonne bonum semen seminasti in agro tuo? Unde ergo habet zizania?".
MATT|13|28|Et ait illis: "Inimicus homo hoc fecit". Servi autem dicunt ei: "Vis, imus et colligimus ea?".
MATT|13|29|Et ait: "Non; ne forte colligentes zizania eradicetis simul cum eis triticum,
MATT|13|30|sinite utraque crescere usque ad messem. Et in tempore messis dicam messoribus: Colligite primum zizania et alligate ea in fasciculos ad comburendum ea, triticum autem congregate in horreum meum" ".
MATT|13|31|Aliam parabolam proposuit eis dicens: " Simile est regnum caelorum grano sinapis, quod accipiens homo seminavit in agro suo.
MATT|13|32|Quod minimum quidem est omnibus seminibus; cum autem creverit, maius est holeribus et fit arbor, ita ut volucres caeli veniant et habitent in ramis eius ".
MATT|13|33|Aliam parabolam locutus est eis: " Simile est regnum caelorum fermento, quod acceptum mulier abscondit in farinae satis tribus, donec fermentatum est totum ".
MATT|13|34|Haec omnia locutus est Iesus in parabolis ad turbas; et sine parabola nihil loquebatur eis,
MATT|13|35|ut adimpleretur, quod dictum erat per prophetam dicentem: Aperiam in parabolis os meum,eructabo abscondita a constitutione mundi ".
MATT|13|36|Tunc, dimissis turbis, venit in domum, et accesserunt ad eum discipuli eius dicentes: " Dissere nobis parabolam zizaniorum agri ".
MATT|13|37|Qui respondens ait: " Qui seminat bonum semen, est Filius hominis;
MATT|13|38|ager autem est mundus; bonum vero semen, hi sunt filii regni; zizania autem filii sunt Mali;
MATT|13|39|inimicus autem, qui seminavit ea, est Diabolus; messis vero consummatio saeculi est; messores autem angeli sunt.
MATT|13|40|Sicut ergo colliguntur zizania et igni comburuntur, sic erit in consummatione saeculi:
MATT|13|41|mittet Filius hominis angelos suos, et colligent de regno eius omnia scandala et eos, qui faciunt iniquitatem,
MATT|13|42|et mittent eos in caminum ignis; ibi erit fletus et stridor dentium.
MATT|13|43|Tunc iusti fulgebunt sicut sol in regno Pa tris eorum. Qui habet aures, audiat.
MATT|13|44|Simile est regnum caelorum thesauro abscondito in agro; quem qui invenit homo abscondit et prae gaudio illius vadit et vendit universa, quae habet, et emit agrum illum.
MATT|13|45|Iterum simile est regnum caelorum homini negotiatori quaerenti bonas margaritas.
MATT|13|46|Inventa autem una pretiosa margarita, abiit et vendidit omnia, quae habuit, et emit eam.
MATT|13|47|Iterum simile est regnum caelorum sagenae missae in mare et ex omni genere congreganti;
MATT|13|48|quam, cum impleta esset, educentes secus litus et sedentes collegerunt bonos in vasa, malos autem foras miserunt.
MATT|13|49|Sic erit in consummatione saeculi: exibunt angeli et separabunt malos de medio iustorum
MATT|13|50|et mittent eos in caminum ignis; ibi erit fletus et stridor dentium.
MATT|13|51|Intellexistis haec omnia? ". Dicunt ei: " Etiam ".
MATT|13|52|Ait autem illis: " Ideo omnis scriba doctus in regno caelorum similis est homini patri familias, qui profert de thesauro suo nova et vetera ".
MATT|13|53|Et factum est, cum consummasset Iesus parabolas istas, transiit inde.
MATT|13|54|Et veniens in patriam suam, docebat eos in synagoga eorum, ita ut mirarentur et dicerent: " Unde huic sapientia haec et virtutes?
MATT|13|55|Nonne hic est fabri filius? Nonne mater eius dicitur Maria, et fratres eius Iacobus et Ioseph et Simon et Iudas?
MATT|13|56|Et sorores eius nonne omnes apud nos sunt? Unde ergo huic omnia ista?.
MATT|13|57|Et scandalizabantur in eo. Iesus autem dixit eis: " Non est propheta sine honore nisi in patria et in domo sua ".
MATT|13|58|Et non fecit ibi virtutes multas propter incredulitatem illorum.
MATT|14|1|In illo tempore audivit He rodes tetrarcha famam Iesu
MATT|14|2|et ait pueris suis: " Hic est Ioannes Baptista; ipse surrexit a mortuis, et ideo virtutes operantur in eo ".
MATT|14|3|Herodes enim tenuit Ioannem et alligavit eum et posuit in carcere propter Herodiadem uxorem Philippi fratris sui.
MATT|14|4|Dicebat enim illi Ioannes: " Non licet tibi habere eam ".
MATT|14|5|Et volens illum occidere, timuit populum, quia sicut prophetam eum habebant.
MATT|14|6|Die autem natalis Herodis saltavit filia Herodiadis in medio et placuit Herodi,
MATT|14|7|unde cum iuramento pollicitus est ei dare, quodcumque postulasset.
MATT|14|8|At illa, praemonita a matre sua: " Da mihi, inquit, hic in disco caput Ioannis Baptistae ".
MATT|14|9|Et contristatus rex propter iuramentum et eos, qui pariter recumbebant, iussit dari
MATT|14|10|misitque et decollavit Ioannem in carcere;
MATT|14|11|et allatum est caput eius in disco et datum est puellae, et tulit matri suae.
MATT|14|12|Et accedentes discipuli eius tulerunt corpus et sepelierunt illud et venientes nuntiaverunt Iesu.
MATT|14|13|Quod cum audisset Iesus, secessit inde in navicula in locum desertum seorsum; et cum audissent, turbae secutae sunt eum pedestres de civitatibus.
MATT|14|14|Et exiens vidit turbam multam et misertus est eorum et curavit languidos eorum.
MATT|14|15|Vespere autem facto, accesserunt ad eum discipuli dicentes: " Desertus est locus, et hora iam praeteriit; dimitte turbas, ut euntes in castella emant sibi escas ".
MATT|14|16|Iesus autem dixit eis: " Non habent necesse ire; date illis vos manducare ".
MATT|14|17|Illi autem dicunt ei: " Non habemus hic nisi quinque panes et duos pisces ".
MATT|14|18|Qui ait: " Afferte illos mihi huc ".
MATT|14|19|Et cum iussisset turbas discumbere supra fenum, acceptis quinque panibus et duobus piscibus, aspiciens in caelum benedixit et fregit et dedit discipulis panes, discipuli autem turbis.
MATT|14|20|Et manducaverunt omnes et saturati sunt; et tulerunt reliquias fragmentorum duodecim cophinos plenos.
MATT|14|21|Manducantium autem fuit numerus fere quinque milia virorum, exceptis mulieribus et parvulis.
MATT|14|22|Et statim iussit discipulos ascendere in naviculam et praecedere eum trans fretum, donec dimitteret turbas.
MATT|14|23|Et dimissis turbis, ascendit in montem solus orare. Vespere autem facto, solus erat ibi.
MATT|14|24|Navicula autem iam multis stadiis a terra distabat, fluctibus iactata; erat enim contrarius ventus.
MATT|14|25|Quarta autem vigilia noctis venit ad eos ambulans supra mare.
MATT|14|26|Discipuli autem, videntes eum supra mare ambulantem, turbati sunt dicentes: " Phantasma est ", et prae timore clamaverunt.
MATT|14|27|Statimque Iesus locutus est eis dicens: " Habete fiduciam, ego sum; nolite timere! ".
MATT|14|28|Respondens autem ei Petrus dixit: " Domine, si tu es, iube me venire ad te super aquas ".
MATT|14|29|At ipse ait: " Veni! ". Et descendens Petrus de navicula ambulavit super aquas et venit ad Iesum.
MATT|14|30|Videns vero ventum validum timuit et, cum coepisset mergi, clamavit dicens: " Domine, salvum me fac! ".
MATT|14|31|Continuo autem Iesus extendens manum apprehendit eum et ait illi: " Modicae fidei, quare dubitasti? ".
MATT|14|32|Et cum ascendissent in naviculam, cessavit ventus.
MATT|14|33|Qui autem in navicula erant, adoraverunt eum dicentes: " Vere Filius Dei es! ".
MATT|14|34|Et cum transfretassent, venerunt in terram Gennesaret.
MATT|14|35|Et cum cognovissent eum viri loci illius, miserunt in universam regionem illam et obtulerunt ei omnes male habentes,
MATT|14|36|et rogabant eum, ut vel fimbriam vestimenti eius tangerent; et, quicumque tetigerunt, salvi facti sunt.
MATT|15|1|Tunc accedunt ad Iesum ab Hierosolymis pharisaei et scribae dicentes:
MATT|15|2|" Quare discipuli tui transgrediuntur traditionem seniorum? Non enim lavant manus suas, cum panem manducant ".
MATT|15|3|Ipse autem respondens ait illis: " Quare et vos transgredimini mandatum Dei propter traditionem vestram?
MATT|15|4|Nam Deus dixit: "Honora patrem tuum et matrem" et: "Qui maledixerit patri vel matri, morte moriatur".
MATT|15|5|Vos autem dicitis: "Quicumque dixerit patri vel matri: Munus est, quodcumque ex me profuerit,
MATT|15|6|non honorificabit patrem suum"; et irritum fecistis verbum Dei propter traditionem vestram.
MATT|15|7|Hypocritae! Bene prophetavit de vobis Isaias dicens:
MATT|15|8|"Populus hic labiis me honorat,cor autem eorum longe est a me;
MATT|15|9|sine causa autem colunt medocentes doctrinas mandata homi num" ".
MATT|15|10|Et convocata ad se turba, dixit eis: " Audite et intellegite:
MATT|15|11|Non quod intrat in os, coinquinat hominem; sed quod procedit ex ore, hoc coinquinat hominem! ".
MATT|15|12|Tunc accedentes discipuli dicunt ei: " Scis quia pharisaei, audito verbo, scandalizati sunt? ".
MATT|15|13|At ille respondens ait: " Omnis plantatio, quam non plantavit Pater meus caelestis, eradicabitur.
MATT|15|14|Sinite illos: caeci sunt, duces caecorum. Caecus autem si caeco ducatum praestet, ambo in foveam cadent ".
MATT|15|15|Respondens autem Petrus dixit ei: " Edissere nobis parabolam istam ".
MATT|15|16|At ille dixit: " Adhuc et vos sine intellectu estis?
MATT|15|17|Non intellegitis quia omne quod in os intrat, in ventrem vadit et in secessum emittitur?
MATT|15|18|Quae autem procedunt de ore, de corde exeunt, et ea coinquinant hominem.
MATT|15|19|De corde enim exeunt cogitationes malae, homicidia, adulteria, fornicationes, furta, falsa testimonia, blasphemiae.
MATT|15|20|Haec sunt, quae coinquinant hominem; non lotis autem manibus manducare non coinquinat hominem ".
MATT|15|21|Et egressus inde Iesus, secessit in partes Tyri et Sidonis.
MATT|15|22|Et ecce mulier Chananaea a finibus illis egressa clamavit dicens: " Miserere mei, Domine, fili David! Filia mea male a daemonio vexatur ".
MATT|15|23|Qui non respondit ei verbum.Et accedentes discipuli eius rogabant eum dicentes: " Dimitte eam, quia clamat post nos ".
MATT|15|24|Ipse autem respondens ait: " Non sum missus nisi ad oves, quae perierunt domus Israel ".
MATT|15|25|At illa venit et adoravit eum dicens: " Domine, adiuva me! ".
MATT|15|26|Qui respondens ait: " Non est bonum sumere panem filiorum et mittere catellis ".
MATT|15|27|At illa dixit: " Etiam, Domine, nam et catelli edunt de micis, quae cadunt de mensa dominorum suorum ".
MATT|15|28|Tunc respondens Iesus ait illi: " O mulier, magna est fides tua! Fiat tibi, sicut vis ". Et sanata est filia illius ex illa hora.
MATT|15|29|Et cum transisset inde, Iesus venit secus mare Galilaeae et ascendens in montem sedebat ibi.
MATT|15|30|Et accesserunt ad eum turbae multae habentes secum claudos, caecos, debiles, mutos et alios multos et proiecerunt eos ad pedes eius, et curavit eos,
MATT|15|31|ita ut turba miraretur videntes mutos loquentes, debiles sanos et claudos ambulantes et caecos videntes. Et magnificabant Deum Israel.
MATT|15|32|Iesus autem convocatis discipulis suis dixit: " Misereor turbae, quia triduo iam perseverant mecum et non habent, quod manducent; et dimittere eos ieiunos nolo, ne forte deficiant in via ".
MATT|15|33|Et dicunt ei discipuli: " Unde nobis in deserto panes tantos, ut saturemus turbam tantam? ".
MATT|15|34|Et ait illis Iesus: " Quot panes habetis? ". At illi dixerunt: " Septem et paucos pisciculos ".
MATT|15|35|Et praecepit turbae, ut discumberet super terram;
MATT|15|36|et accipiens septem panes et pisces et gratias agens fregit et dedit discipulis, discipuli autem turbis.
MATT|15|37|Et comederunt omnes et saturati sunt; et, quod superfuit de fragmentis, tulerunt septem sportas plenas.
MATT|15|38|Erant autem, qui manducaverant, quattuor milia hominum extra mulieres et parvulos.
MATT|15|39|Et dimissis turbis, ascendit in naviculam et venit in fines Magadan.
MATT|16|1|Et accesserunt ad eum pharisaei et sadducaei tentantes et rogaverunt eum, ut signum de caelo ostenderet eis.
MATT|16|2|At ille respondens ait eis: " Facto vespere dicitis: "Serenum erit, rubicundum est enim caelum";
MATT|16|3|et mane: "Hodie tempestas, rutilat enim triste caelum". Faciem quidem caeli diiudicare nostis, signa autem temporum non potestis.
MATT|16|4|Generatio mala et adultera signum quaerit, et signum non dabitur ei, nisi signum Ionae ". Et, relictis illis, abiit.
MATT|16|5|Et cum venissent discipuli trans fretum, obliti sunt panes accipere.
MATT|16|6|Iesus autem dixit illis: " Intuemini et cavete a fermento pharisaeorum et sadducaeorum ".
MATT|16|7|At illi cogitabant inter se dicentes: " Panes non accepimus!".
MATT|16|8|Sciens autem Iesus dixit: " Quid cogitatis inter vos, modicae fidei, quia panes non habetis?
MATT|16|9|Nondum intellegitis neque recordamini quinque panum quinque milium hominum, et quot cophinos sumpsistis?
MATT|16|10|Neque septem panum quattuor milium hominum, et quot sportas sumpsistis?
MATT|16|11|Quomodo non intellegitis quia non de panibus dixi vobis? Sed cavete a fermento pharisaeorum et sadducaeorum ".
MATT|16|12|Tunc intellexerunt quia non dixerit cavendum a fermento panum sed a doctrina pharisaeorum et sadducaeorum.
MATT|16|13|Venit autem Iesus in partes Caesareae Philippi et interrogabat discipulos suos dicens: " Quem dicunt homines esse Filium hominis?".
MATT|16|14|At illi dixerunt: " Alii Ioannem Baptistam, alii autem Eliam, alii vero Ieremiam, aut unum ex prophetis ".
MATT|16|15|Dicit illis: " Vos autem quem me esse dicitis? ".
MATT|16|16|Respondens Simon Petrus dixit: " Tu es Christus, Filius Dei vivi ".
MATT|16|17|Respondens autem Iesus dixit ei: " Beatus es, Simon Bariona, quia caro et sanguis non revelavit tibi sed Pater meus, qui in caelis est.
MATT|16|18|Et ego dico tibi: Tu es Petrus, et super hanc petram aedificabo Ecclesiam meam; et portae inferi non praevalebunt adversum eam.
MATT|16|19|Tibi dabo claves regni caelorum; et quodcumque ligaveris super terram, erit ligatum in caelis, et quodcumque solveris super terram, erit solutum in caelis ".
MATT|16|20|Tunc praecepit discipulis, ut nemini dicerent quia ipse esset Christus.
MATT|16|21|Exinde coepit Iesus ostendere discipulis suis quia oporteret eum ire Hierosolymam et multa pati a senioribus et principibus sacerdotum et scribis et occidi et tertia die resurgere.
MATT|16|22|Et assumens eum Petrus coepit increpare illum dicens: " Absit a te, Domine; non erit tibi hoc ".
MATT|16|23|Qui conversus dixit Petro: " Vade post me, Satana! Scandalum es mihi, quia non sapis ea, quae Dei sunt, sed ea, quae hominum! ".
MATT|16|24|Tunc Iesus dixit discipulis suis: " Si quis vult post me venire, abneget semetipsum et tollat crucem suam et sequatur me.
MATT|16|25|Qui enim voluerit animam suam salvam facere, perdet eam; qui autem perdiderit animam suam propter me, inveniet eam.
MATT|16|26|Quid enim prodest homini, si mundum universum lucretur, animae vero suae detrimentum patiatur? Aut quam dabit homo commutationem pro anima sua?
MATT|16|27|Filius enim hominis venturus est in gloria Patris sui cum angelis suis, et tunc reddet unicuique secundum opus eius.
MATT|16|28|Amen dico vobis: Sunt quidam de hic stantibus, qui non gustabunt mortem, donec videant Filium hominis venientem in regno suo ".
MATT|17|1|Et post dies sex assumit Iesus Petrum et Iacobum et Ioan nem fratrem eius et ducit illos in montem excelsum seorsum.
MATT|17|2|Et transfiguratus est ante eos; et resplenduit facies eius sicut sol, vestimenta autem eius facta sunt alba sicut lux.
MATT|17|3|Et ecce apparuit illis Moyses et Elias cum eo loquentes.
MATT|17|4|Respondens autem Petrus dixit ad Iesum: " Domine, bonum est nos hic esse. Si vis, faciam hic tria tabernacula: tibi unum et Moysi unum et Eliae unum ".
MATT|17|5|Adhuc eo loquente, ecce nubes lucida obumbravit eos; et ecce vox de nube dicens: " Hic est Filius meus dilectus, in quo mihi bene complacui; ipsum audite ".
MATT|17|6|Et audientes discipuli ceciderunt in faciem suam et timuerunt valde.
MATT|17|7|Et accessit Iesus et tetigit eos dixitque eis: " Surgite et nolite timere ".
MATT|17|8|Levantes autem oculos suos, neminem viderunt nisi solum Iesum.
MATT|17|9|Et descendentibus illis de monte, praecepit eis Iesus dicens: " Nemini dixeritis visionem, donec Filius hominis a mortuis resurgat ".
MATT|17|10|Et interrogaverunt eum discipuli dicentes: " Quid ergo scribae dicunt quod Eliam oporteat primum venire? ".
MATT|17|11|At ille respondens ait: " Elias quidem venturus est et restituet omnia.
MATT|17|12|Dico autem vobis quia Elias iam venit, et non cognoverunt eum, sed fecerunt in eo, quaecumque voluerunt; sic et Filius hominis passurus est ab eis ".
MATT|17|13|Tunc intellexerunt discipuli quia de Ioanne Baptista dixisset eis.
MATT|17|14|Et cum venissent ad turbam, accessit ad eum homo genibus provolutus ante eum
MATT|17|15|et dicens: " Domine, miserere filii mei, quia lunaticus est et male patitur; nam saepe cadit in ignem et crebro in aquam.
MATT|17|16|Et obtuli eum discipulis tuis, et non potuerunt curare eum ".
MATT|17|17|Respondens autem Iesus ait: " O generatio incredula et perversa, quousque ero vobiscum? Usquequo patiar vos? Afferte huc illum ad me ".
MATT|17|18|Et increpavit eum Iesus, et exiit ab eo daemonium, et curatus est puer ex illa hora.
MATT|17|19|Tunc accesserunt discipuli ad Iesum secreto et dixerunt: " Quare nos non potuimus eicere illum? ".
MATT|17|20|Ille autem dicit illis: " Propter modicam fidem vestram. Amen quippe dico vobis: Si habueritis fidem sicutgranum sinapis, dicetis monti huic: "Transi hinc illuc!", et transibit, et nihil impossibile erit vobis ".
MATT|17|21|()
MATT|17|22|Conversantibus autem eis in Galilaea, dixit illis Iesus: " Filius hominis tradendus est in manus hominum,
MATT|17|23|et occident eum, et tertio die resurget ". Et contristati sunt vehementer.
MATT|17|24|Et cum venissent Capharnaum, accesserunt, qui didrachma accipiebant, ad Petrum et dixerunt: " Magister vester non solvit didrachma? ".
MATT|17|25|Ait: " Etiam". Et cum intrasset domum, praevenit eum Iesus dicens: " Quid tibi videtur, Simon? Reges terrae a quibus accipiunt tributum vel censum? A filiis suis an ab alienis? ".
MATT|17|26|Cum autem ille dixisset: " Ab alienis ", dixit illi Iesus: " Ergo liberi sunt filii.
MATT|17|27|Ut autem non scandalizemus eos, vade ad mare et mitte hamum; et eum piscem, qui primus ascenderit, tolle; et, aperto ore, eius invenies staterem. Illum sumens, da eis pro me et te ".
MATT|18|1|In illa hora accesserunt di scipuli ad Iesum dicentes: " Quis putas maior est in regno caelorum? ".
MATT|18|2|Et advocans parvulum, statuit eum in medio eorum
MATT|18|3|et dixit: " Amen dico vobis: Nisi conversi fueritis et efiiciamini sicut parvuli, non intrabitis in regnum caelorum.
MATT|18|4|Quicumque ergo humiliaverit se sicut parvulus iste, hic est maior in regno caelorum.
MATT|18|5|Et, qui susceperit unum parvulum talem in nomine meo, me suscipit.
MATT|18|6|Qui autem scandalizaverit unum de pusillis istis, qui in me credunt, expedit ei, ut suspendatur mola asinaria in collo eius et demergatur in profundum maris.
MATT|18|7|Vae mundo ab scandalis! Necesse est enim ut veniant scandala; verumtamen vae homini, per quem scandalum venit!
MATT|18|8|Si autem manus tua vel pes tuus scandalizat te, abscide eum et proice abs te: bonum tibi est ad vitam ingredi debilem vel claudum, quam duas manus vel duos pedes habentem mitti in ignem aeternum.
MATT|18|9|Et si oculus tuus scandalizat te, erue eum et proice abs te: bonum tibi est unoculum in vitam intrare, quam duos oculos habentem mitti in gehennam ignis.
MATT|18|10|Videte, ne contemnatis unum ex his pusillis; dico enim vobis quia angeli eorum in caelis sempervident faciem Patris mei, qui in caelis est.
MATT|18|11|()
MATT|18|12|Quid vobis videtur? Si fuerint alicui centum oves, et erraverit una ex eis, nonne relinquet nonaginta novem in montibus et vadit quaerere eam, quae erravit?
MATT|18|13|Et si contigerit ut inveniat eam, amen dico vobis quia gaudebit super eam magis quam super nonaginta novem, quae non erraverunt.
MATT|18|14|Sic non est voluntas ante Patrem vestrum, qui in caelis est, ut pereat unus de pusillis istis.
MATT|18|15|Si autem peccaverit in te frater tuus, vade, corripe eum inter te et ipsum solum. Si te audierit, lucratus es fratrem tuum;
MATT|18|16|si autem non audierit, adhibe tecum adhuc unum vel duos, ut in ore duorum testium vel trium stet omne verbum;
MATT|18|17|quod si noluerit audire eos, dic ecclesiae; si autem et ecclesiam noluerit audire, sit tibi sicut ethnicus et publicanus.
MATT|18|18|Amen dico vobis: Quaecumque alligaveritis super terram, erunt ligata in caelo; et, quaecumque solveritis super terram, erunt soluta in caelo.
MATT|18|19|Iterum dico vobis: Si duo ex vobis consenserint super terram de omni re, quamcumque petierint, fiet illis a Patre meo, qui in caelis est.
MATT|18|20|Ubi enim sunt duo vel tres congregati in nomine meo, ibi sum in medio eorum ".
MATT|18|21|Tunc accedens Petrus dixit ei: " Domine, quotiens peccabit in me frater meus, et dimittam ei? Usque septies? ".
MATT|18|22|Dicit illi Iesus: " Non dico tibi usque septies sed usque septuagies septies.
MATT|18|23|Ideo assimilatum est regnum caelorum homini regi, qui voluit rationem ponere cum servis suis.
MATT|18|24|Et cum coepisset rationem ponere, oblatus est ei unus, qui debebat decem milia talenta.
MATT|18|25|Cum autem non haberet, unde redderet, iussit eum dominus venumdari et uxorem et filios et omnia, quae habebat, et reddi.
MATT|18|26|Procidens igitur servus ille adorabat eum dicens: "Patientiam habe in me, et omnia reddam tibi".
MATT|18|27|Misertus autem dominus servi illius dimisit eum et debitum dimisit ei.
MATT|18|28|Egressus autem servus ille invenit unum de conservis suis, qui debebat ei centum denarios, et tenens suffocabat eum dicens: "Redde, quod debes!".
MATT|18|29|Procidens igitur conservus eius rogabat eum dicens: "Patientiam habe in me, et reddam tibi".
MATT|18|30|Ille autem noluit, sed abiit et misit eum in carcerem, donec redderet debitum.
MATT|18|31|Videntes autem conservi eius, quae fiebant, contristati sunt valde et venerunt et narraverunt domino suo omnia, quae facta erant.
MATT|18|32|Tunc vocavit illum dominus suus et ait illi: "Serve nequam, omne debitum illud dimisi tibi, quoniam rogasti me;
MATT|18|33|non oportuit et te misereri conservi tui, sicut et ego tui misertus sum?".
MATT|18|34|Et iratus dominus eius tradidit eum tortoribus, quoadusque redderet universum debitum.
MATT|18|35|Sic et Pater meus caelestis faciet vobis, si non remiseritis unusquisque fratri suo de cordibus vestris ".
MATT|19|1|Et factum est, cum consum masset Iesus sermones istos, migravit a Galilaea et venit in fines Iudaeae trans Iordanem.
MATT|19|2|Et secutae sunt eum turbae multae, et curavit eos ibi.
MATT|19|3|Et accesserunt ad eum pharisaei tentantes eum et dicentes: " Licet homini dimittere uxorem suam quacumque ex causa? ".
MATT|19|4|Qui respondens ait: " Non legistis quia, qui creavit ab initio, masculum et feminam fecit eos
MATT|19|5|et dixit: "Propter hoc dimittet homo patrem et matrem et adhaerebit uxori suae, et erunt duo in carne una?".
MATT|19|6|Itaque iam non sunt duo sed una caro. Quod ergo Deus coniunxit, homo non separet ".
MATT|19|7|Dicunt illi: " Quid ergo Moyses mandavit dari libellum repudii et dimittere? ".
MATT|19|8|Ait illis: " Moyses ad duritiam cordis vestri permisit vobis dimittere uxores vestras; ab initio autem non sic fuit.
MATT|19|9|Dico autem vobis quia quicumque dimiserit uxorem suam, nisi ob fornicationem, et aliam duxerit, moechatur ".
MATT|19|10|Dicunt ei discipuli eius: " Si ita est causa hominis cum uxore, non expedit nubere ".
MATT|19|11|Qui dixit eis: " Non omnes capiunt verbum istud, sed quibus datum est.
MATT|19|12|Sunt enim eunuchi, qui de matris utero sic nati sunt; et sunt eunuchi, qui facti sunt ab hominibus; et sunt eunuchi, qui seipsos castraverunt propter regnum caelorum. Qui potest capere, capiat ".
MATT|19|13|Tunc oblati sunt ei parvuli, ut manus eis imponeret et oraret; discipuli autem increpabant eis.
MATT|19|14|Iesus vero ait: " Sinite parvulos et nolite eos prohibere ad me venire; talium est enim regnum caelorum ".
MATT|19|15|Et cum imposuisset eis manus, abiit inde.
MATT|19|16|Et ecce unus accedens ait illi: " Magister, quid boni faciam, ut habeam vitam aeternam? ". Qui dixit ei:
MATT|19|17|" Quid me interrogas de bono? Unus est bonus. Si autem vis ad vitam ingredi, serva mandata ".
MATT|19|18|Dicit illi: " Quae? ". Iesus autem dixit: " Non homicidium facies, non adulterabis, non facies furtum, non falsum testimonium dices,
MATT|19|19|honora patrem et matrem et diliges proximum tuum sicut teipsum ".
MATT|19|20|Dicit illi adulescens: " Omnia haec custodivi. Quid adhuc mihi deest?.
MATT|19|21|Ait illi Iesus: " Si vis perfectus esse, vade, vende, quae habes, et da pauperibus, et habebis thesaurum in caelo; et veni, sequere me ".
MATT|19|22|Cum audisset autem adulescens verbum, abiit tristis; erat enim habens multas possessiones.
MATT|19|23|Iesus autem dixit discipulis suis: " Amen dico vobis: Dives difficile intrabit in regnum caelorum.
MATT|19|24|Et iterum dico vobis: Facilius est camelum per foramen acus transire, quam divitem intrare in regnum Dei ".
MATT|19|25|Auditis autem his, discipuli mirabantur valde dicentes: " Quis ergo poterit salvus esse? ".
MATT|19|26|Aspiciens autem Iesus dixit illis: " Apud homines hoc impossibile est, apud Deum autem omnia possibilia sunt ".
MATT|19|27|Tunc respondens Petrus dixit ei: " Ecce nos reliquimus omnia et secuti sumus te. Quid ergo erit nobis? ".
MATT|19|28|Iesus autem dixit illis: " Amen dico vobis quod vos, qui secuti estis me, in regeneratione, cum sederit Filius hominis in throno gloriae suae, sedebitis et vos super thronos duodecim, iudicantes duodecim tribus Israel.
MATT|19|29|Et omnis, qui reliquit domos vel fratres aut sorores aut patrem aut matrem aut filios aut agros propter nomen meum, centuplum accipiet et vitam aeternam possidebit.
MATT|19|30|Multi autem erunt primi novissimi, et novissimi primi.
MATT|20|1|Simile est enim regnum cae lorum homini patri familias, qui exiit primo mane conducere operarios in vineam suam;
MATT|20|2|conventione autem facta cum operariis ex denario diurno, misit eos in vineam suam.
MATT|20|3|Et egressus circa horam tertiam vidit alios stantes in foro otiosos
MATT|20|4|et illis dixit: "Ite et vos in vineam; et, quod iustum fuerit, dabo vobis".
MATT|20|5|Illi autem abierunt. Iterum autem exiit circa sextam et nonam horam et fecit similiter.
MATT|20|6|Circa undecimam vero exiit et invenit alios stantes et dicit illis: Quid hic statis tota die otiosi?".
MATT|20|7|Dicunt ei: "Quia nemo nos conduxit". Dicit illis: "Ite et vos in vineam".
MATT|20|8|Cum sero autem factum esset, dicit dominus vineae procuratori suo: " Voca operarios et redde illis mercedem incipiens a novissimis usque ad primos ".
MATT|20|9|Et cum venissent, qui circa undecimam horam venerant, acceperunt singuli denarium.
MATT|20|10|Venientes autem primi arbitrati sunt quod plus essent accepturi; acceperunt autem et ipsi singuli denarium.
MATT|20|11|Accipientes autem murmurabant adversus patrem familias
MATT|20|12|dicentes: "Hi novissimi una hora fecerunt, et pares illos nobis fecisti, qui portavimus pondus diei et aestum!".
MATT|20|13|At ille respondens uni eorum dixit: "Amice, non facio tibi iniuriam; nonne ex denario convenisti mecum?
MATT|20|14|Tolle, quod tuum est, et vade; volo autem et huic novissimo dare sicut et tibi.
MATT|20|15|Aut non licet mihi, quod volo, facere de meis? An oculus tuus nequam est, quia ego bonus sum?".
MATT|20|16|Sic erunt novissimi primi, et primi novissimi ".
MATT|20|17|Et ascendens Iesus Hierosolymam assumpsit Duodecim discipulos secreto et ait illis in via:
MATT|20|18|" Ecce ascendimus Hierosolymam, et Filius hominis tradetur principibus sacerdotum et scribis, et condemnabunt eum morte
MATT|20|19|et tradent eum gentibus ad illudendum et flagellandum et crucifigendum, et tertia die resurget ".
MATT|20|20|Tunc accessit ad eum mater filiorum Zebedaei cum filiis suis, adorans et petens aliquid ab eo.
MATT|20|21|Qui dixit ei: " Quid vis? ". Ait illi: " Dic ut sedeant hi duo filii mei unus ad dexteram tuam et unus ad sinistram in regno tuo ".
MATT|20|22|Respondens autem Iesus dixit: " Nescitis quid petatis. Potestis bibere calicem, quem ego bibiturus sum? ". Dicunt ei: " Possumus ".
MATT|20|23|Ait illis: " Calicem quidem meum bibetis, sedere autem ad dexteram meam et sinistram non est meum dare illud, sed quibus paratum est a Patre meo.
MATT|20|24|Et audientes decem indignati sunt de duobus fratribus.
MATT|20|25|Iesus autem vocavit eos ad se et ait: " Scitis quia principes gentium dominantur eorum et, qui magni sunt, potestatem exercent in eos.
MATT|20|26|Non ita erit inter vos, sed quicumque voluerit inter vos magnus fieri, erit vester minister;
MATT|20|27|et, quicumque voluerit inter vos primus esse, erit vester servus;
MATT|20|28|sicut Filius hominis non venit ministrari sed ministrare et dare animam suam redemptionem pro multis ".
MATT|20|29|Et egredientibus illis ab Iericho, secuta est eum turba multa.
MATT|20|30|Et ecce duo caeci sedentes secus viam audierunt quia Iesus transiret et clamaverunt dicentes: " Domine, miserere nostri, fili David! ".
MATT|20|31|Turba autem increpabat eos, ut tacerent; at illi magis clamabant dicentes: " Domine, miserere nostri, fili David! ".
MATT|20|32|Et stetit Iesus et vocavit eos et ait: " Quid vultis, ut faciam vobis?".
MATT|20|33|Dicunt illi: " Domine, ut aperiantur oculi nostri ".
MATT|20|34|Misertus autem Iesus, tetigit oculos eorum; et confestim viderunt et secuti sunt eum.
MATT|21|1|Et cum appropinquassent Hierosolymis et venissent Bethfage, ad montem Oliveti, tunc Iesus misit duos discipulos
MATT|21|2|dicens eis: " Ite in castellum, quod contra vos est, et statim invenietis asinam alligatam et pullum cum ea; solvite et adducite mihi.
MATT|21|3|Et si quis vobis aliquid dixerit, dicite: "Dominus eos necessarios habet", et confestim dimittet eos ".
MATT|21|4|Hoc autem factum est, ut impleretur, quod dictum est per prophetam dicentem:
MATT|21|5|" Dicite filiae Sion:Ecce Rex tuus venit tibi,mansuetus et sedens super asinamet super pullum filium subiugalis ".
MATT|21|6|Euntes autem discipuli fecerunt, sicut praecepit illis Iesus,
MATT|21|7|et adduxerunt asinam et pullum; et imposuerunt super eis vestimenta sua, et sedit super ea.
MATT|21|8|Plurima autem turba straverunt vestimenta sua in via; alii autem caedebant ramos de arboribus et sternebant in via.
MATT|21|9|Turbae autem, quae praecedebant eum et quae sequebantur, clamabant dicentes: " Hosanna filio David! Benedictus, qui venit in nomine Domini! Hosanna in altissimis! ".
MATT|21|10|Et cum intrasset Hierosolymam, commota est universa civitas dicens: " Quis est hic?".
MATT|21|11|Turbae autem dicebant: " Hic est Iesus propheta a Nazareth Galilaeae ".
MATT|21|12|Et intravit Iesus in templum et eiciebat omnes vendentes et ementes in templo, et mensas nummulariorum evertit et cathedras vendentium columbas,
MATT|21|13|et dicit eis: " Scriptum est: "Domus mea domus orationis vocabitur". Vos autem facitis eam speluncam latronum ".
MATT|21|14|Et accesserunt ad eum caeci et claudi in templo, et sanavit eos.
MATT|21|15|Videntes autem principes sacerdotum et scribae mirabilia, quae fecit, et pueros clamantes in templo et dicentes: " Hosanna filio David ", indignati sunt
MATT|21|16|et dixerunt ei: " Audis quid isti dicant? ". Iesus autem dicit eis: " Utique; numquam legistis: "Ex ore infantium et lactantium perfecisti laudem"? ".
MATT|21|17|Et relictis illis, abiit foras extra civitatem in Bethaniam ibique mansit.
MATT|21|18|Mane autem revertens in civitatem, esuriit.
MATT|21|19|Et videns fici arborem unam secus viam, venit ad eam; et nihil invenit in ea nisi folia tantum et ait illi: " Numquam ex te fructus nascatur in sempiternum ". Et arefacta est continuo ficulnea.
MATT|21|20|Et videntes discipuli mirati sunt dicentes: " Quomodo continuo aruit ficulnea? ".
MATT|21|21|Respondens autem Iesus ait eis: " Amen dico vobis: Si habueritis fidem et non haesitaveritis, non solum de ficulnea facietis, sed et si monti huic dixeritis: "Tolle et iacta te in mare", fiet.
MATT|21|22|Et omnia, quaecumque petieritis in oratione credentes, accipietis ".
MATT|21|23|Et cum venisset in templum, accesserunt ad eum docentem principes sacerdotum et seniores populi dicentes: " In qua potestate haec facis? Et quis tibi dedit hanc potestatem? ".
MATT|21|24|Respondens autem Iesus dixit illis: " Interrogabo vos et ego unum sermonem, quem si dixeritis mihi, et ego vobis dicam, in qua potestate haec facio:
MATT|21|25|Baptismum Ioannis unde erat? A caelo an ex hominibus? ". At illi cogitabant inter se dicentes: " Si dixerimus: "E caelo", dicet nobis: Quare ergo non credidistis illi?";
MATT|21|26|si autem dixerimus: "Ex hominibus", timemus turbam; omnes enim habent Ioannem sicut prophetam ".
MATT|21|27|Et respondentes Iesu dixerunt: " Nescimus ". Ait illis et ipse: " Nec ego dico vobis in qua potestate haec facio ".
MATT|21|28|" Quid autem vobis videtur? Homo quidam habebat duos filios. Et accedens ad primum dixit: "Fili, vade hodie, operare in vinea".
MATT|21|29|Ille autem respondens ait: "Nolo"; postea autem paenitentia motus abiit.
MATT|21|30|Accedens autem ad alterum dixit similiter. At ille respondens ait: "Eo, domine"; et non ivit.
MATT|21|31|Quis ex duobus fecit voluntatem patris? ". Dicunt: " Primus ". Dicit illis Iesus: " Amen dico vobis: Publicani et meretrices praecedunt vos in regnum Dei.
MATT|21|32|Venit enim ad vos Ioannes in via iustitiae, et non credidistis ei; publicani autem et meretrices crediderunt ei. Vos autem videntes nec paenitentiam habuistis postea, ut crederetis ei.
MATT|21|33|Aliam parabolam audite. Homo erat pater familias, qui plantavit vineam et saepem circumdedit ei et fodit in ea torcular et aedificavit turrim et locavit eam agricolis et peregre profectus est.
MATT|21|34|Cum autem tempus fructuum appropinquasset, misit servos suos ad agricolas, ut acciperent fructus eius.
MATT|21|35|Et agricolae, apprehensis servis eius, alium ceciderunt, alium occiderunt, alium vero lapidaverunt.
MATT|21|36|Iterum misit alios servos plures prioribus, et fecerunt illis similiter.
MATT|21|37|Novissime autem misit ad eos filium suum dicens: "Verebuntur filium meum".
MATT|21|38|Agricolae autem videntes filium dixerunt intra se: "Hic est heres. Venite, occidamus eum et habebimus hereditatem eius".
MATT|21|39|Et apprehensum eum eiecerunt extra vineam et occiderunt.
MATT|21|40|Cum ergo venerit dominus vineae, quid faciet agricolis illis? ".
MATT|21|41|Aiunt illi: " Malos male perdet et vineam locabit aliis agricolis, qui reddant ei fructum temporibus suis ".
MATT|21|42|Dicit illis Iesus: " Numquam legistis in Scripturis:Lapidem quem reprobaverunt aedificantes,hic factus est in caput anguli;a Domino factum est istudet est mirabile in oculis nostris"?
MATT|21|43|Ideo dico vobis quia auferetur a vobis regnum Dei et dabitur genti facienti fructus eius.
MATT|21|44|Et, qui ceciderit super lapidem istum confringetur; super quem vero ceciderit, conteret eum ".
MATT|21|45|Et cum audissent principes sacerdotum et pharisaei parabolas eius, cognoverunt quod de ipsis diceret;
MATT|21|46|et quaerentes eum tenere, timuerunt turbas, quoniam sicut prophetam eum habebant.
MATT|22|1|Et respondens Iesus dixit ite rum in parabolis eis dicens:
MATT|22|2|" Simile factum est regnum caelorum homini regi, qui fecit nuptias filio suo.
MATT|22|3|Et misit servos suos vocare invitatos ad nuptias, et nolebant venire.
MATT|22|4|Iterum misit alios servos dicens: "Dicite invitatis: Ecce prandium meum paravi, tauri mei et altilia occisa, et omnia parata; venite ad nuptias".
MATT|22|5|Illi autem neglexerunt et abierunt, alius in villam suam, alius vero ad negotiationem suam;
MATT|22|6|reliqui vero tenuerunt servos eius et contumelia affectos occiderunt.
MATT|22|7|Rex autem iratus est et, missis exercitibus suis, perdidit homicidas illos et civitatem illorum succendit.
MATT|22|8|Tunc ait servis suis: "Nuptiae quidem paratae sunt, sed qui invitati erant, non fuerunt digni;
MATT|22|9|ite ergo ad exitus viarum, et quoscumque inveneritis, vocate ad nuptias".
MATT|22|10|Et egressi servi illi in vias, congregaverunt omnes, quos invenerunt, malos et bonos; et impletae sunt nuptiae discumbentium.
MATT|22|11|Intravit autem rex, ut videret discumbentes, et vidit ibi hominem non vestitum veste nuptiali
MATT|22|12|et ait illi: "Amice, quomodo huc intrasti, non habens vestem nuptialem?". At ille obmutuit.
MATT|22|13|Tunc dixit rex ministris: "Ligate pedes eius et manus et mittite eum in tenebras exteriores: ibi erit fletus et stridor dentium".
MATT|22|14|Multi enim sunt vocati, pauci vero electi ".
MATT|22|15|Tunc abeuntes pharisaei consilium inierunt, ut caperent eum in sermone.
MATT|22|16|Et mittunt ei discipulos suos cum herodianis dicentes: " Magister, scimus quia verax es et viam Dei in veritate doces, et non est tibi cura de aliquo; non enim respicis personam hominum.
MATT|22|17|Dic ergo nobis quid tibi videatur: Licet censum dare Caesari an non? ".
MATT|22|18|Cognita autem Iesus nequitia eorum, ait: " Quid me tentatis, hypocritae?
MATT|22|19|Ostendite mihi nomisma census ". At illi obtulerunt ei denarium.
MATT|22|20|Et ait illis: " Cuius est imago haec et suprascriptio? ".
MATT|22|21|Dicunt ei: " Caesaris ". Tunc ait illis: " Reddite ergo, quae sunt Caesaris, Caesari et, quae sunt Dei, Deo ".
MATT|22|22|Et audientes mirati sunt et, relicto eo, abierunt.
MATT|22|23|In illo die accesserunt ad eum sadducaei, qui dicunt non esse resurrectionem, et interrogaverunt eum
MATT|22|24|dicentes: " Magister, Moyses dixit, si quis mortuus fuerit non habens filios, ut ducat frater eius uxorem illius et suscitet semen fratri suo.
MATT|22|25|Erant autem apud nos septem fratres: et primus, uxore ducta, defunctus est et non habens semen reliquit uxorem suam fratri suo;
MATT|22|26|similiter secundus et tertius usque ad septimum.
MATT|22|27|Novissime autem omnium mulier defuncta est.
MATT|22|28|In resurrectione ergo cuius erit de septem uxor? Omnes enim habuerunt eam ".
MATT|22|29|Respondens autem Iesus ait illis: " Erratis nescientes Scripturas neque virtutem Dei;
MATT|22|30|in resurrectione enim neque nubent neque nubentur, sed sunt sicut angeli in caelo.
MATT|22|31|De resurrectione autem mortuorum non legistis, quod dictum est vobis a Deo dicente:
MATT|22|32|"Ego sum Deus Abraham et Deus Isaac et Deus Iacob"? Non est Deus mortuorum sed viventium ".
MATT|22|33|Et audientes turbae mirabantur in doctrina eius.
MATT|22|34|Pharisaei autem audientes quod silentium imposuisset sadducaeis, convenerunt in unum.
MATT|22|35|Et interrogavit unus ex eis legis doctor tentans eum:
MATT|22|36|" Magister, quod est mandatum magnum in Lege? ".
MATT|22|37|Ait autem illi: " Diliges Dominum Deum tuum in toto corde tuo et in tota anima tua et in tota mente tua:
MATT|22|38|hoc est magnum et primum mandatum.
MATT|22|39|Secundum autem simile est huic: Diliges proximum tuum sicut teipsum.
MATT|22|40|In his duobus mandatis universa Lex pendet et Prophetae ".
MATT|22|41|Congregatis autem pharisaeis, interrogavit eos Iesus
MATT|22|42|dicens: " Quid vobis videtur de Christo? Cuius filius est? ". Dicunt ei: " David ".
MATT|22|43|Ait illis: " Quomodo ergo David in Spiritu vocat eum Dominum dicens:
MATT|22|44|"Dixit Dominus Domino meo: Sede a dextris meis,donec ponam inimicos tuos sub pedibus tuis"?
MATT|22|45|Si ergo David vocat eum Dominum, quomodo filius eius est? ".
MATT|22|46|Et nemo poterat respondere ei verbum, neque ausus fuit quisquam ex illa die eum amplius interrogare.
MATT|23|1|Tunc Iesus locutus est ad turbas et ad discipulos suos
MATT|23|2|dicens: " Super cathedram Moysis sederunt scribae et pharisaei.
MATT|23|3|Omnia ergo, quaecumque dixerint vobis, facite et servate; secundum opera vero eorum nolite facere: dicunt enim et non faciunt.
MATT|23|4|Alligant autem onera gravia et importabilia et imponunt in umeros hominum, ipsi autem digito suo nolunt ea movere.
MATT|23|5|Omnia vero opera sua faciunt, ut videantur ab hominibus: dilatant enim phylacteria sua et magnificant fimbrias,
MATT|23|6|amant autem primum recubitum in cenis et primas cathedras in synagogis
MATT|23|7|et salutationes in foro et vocari ab hominibus Rabbi.
MATT|23|8|Vos autem nolite vocari Rabbi; unus enim est Magister vester, omnes autem vos fratres estis.
MATT|23|9|Et Patrem nolite vocare vobis super terram, unus enim est Pater vester, caelestis.
MATT|23|10|Nec vocemini Magistri, quia Magister vester unus est, Christus.
MATT|23|11|Qui maior est vestrum, erit minister vester.
MATT|23|12|Qui autem se exaltaverit, humiliabitur; et, qui se humiliaverit, exaltabitur.
MATT|23|13|Vae autem vobis, scribae et pharisaei hypocritae, quia clauditis regnum caelorum ante homines! Vosenim non intratis nec introeuntes sinitis intrare.
MATT|23|14|()
MATT|23|15|Vae vobis, scribae et pharisaei hypocritae, quia circuitis mare et aridam, ut faciatis unum proselytum, et cum fuerit factus, facitis eum filium gehennae duplo quam vos!
MATT|23|16|Vae vobis, duces caeci, qui dicitis: "Quicumque iuraverit per templum, nihil est; quicumque autem iuraverit in auro templi, debet".
MATT|23|17|Stulti et caeci! Quid enim maius est: aurum an templum, quod sanctificat aurum?
MATT|23|18|Et: "Quicumque iuraverit in altari, nihil est; quicumque autem iuraverit in dono, quod est super illud, debet".
MATT|23|19|Caeci! Quid enim maius est: donum an altare, quod sanctificat donum?
MATT|23|20|Qui ergo iuraverit in altari, iurat in eo et in omnibus, quae super illud sunt;
MATT|23|21|et, qui iuraverit in templo, iurat in illo et in eo, qui inhabitat in ipso;
MATT|23|22|et, qui iuraverit in caelo, iurat in throno Dei et in eo, qui sedet super eum.
MATT|23|23|Vae vobis, scribae et pharisaei hypocritae, quia decimatis mentam et anethum et cyminum et reliquistis, quae graviora sunt legis: iudicium et misericordiam et fidem! Haec oportuit facere et illa non omittere.
MATT|23|24|Duces caeci, excolantes culicem, camelum autem glutientes.
MATT|23|25|Vae vobis, scribae et pharisaei hypocritae, quia mundatis, quod de foris est calicis et paropsidis, intus autem pleni sunt rapina et immunditia!
MATT|23|26|Pharisaee caece, munda prius, quod intus est calicis, ut fiat et id, quod de foris eius est, mundum.
MATT|23|27|Vae vobis, scribae et pharisaei hypocritae, quia similes estis sepulcris dealbatis, quae a foris quidem parent speciosa, intus vero plena sunt ossibus mortuorum et omni spurcitia!
MATT|23|28|Sic et vos a foris quidem paretis hominibus iusti, intus autem pleni estis hypocrisi et iniquitate.
MATT|23|29|Vae vobis, scribae et pharisaei hypocritae, qui aedificatis sepulcra prophetarum et ornatis monumenta iustorum
MATT|23|30|et dicitis: "Si fuissemus in diebus patrum nostrorum, non essemus socii eorum in sanguine prophetarum"!
MATT|23|31|Itaque testimonio estis vobismetipsis quia filii estis eorum, qui prophetas occiderunt.
MATT|23|32|Et vos implete mensuram patrum vestrorum.
MATT|23|33|Serpentes, genimina viperarum, quomodo fugietis a iudicio gehennae?
MATT|23|34|Ideo ecce ego mitto ad vos prophetas et sapientes et scribas; ex illis occidetis et crucifigetis et ex eis flagellabitis in synagogis vestris et persequemini de civitate in civitatem,
MATT|23|35|ut veniat super vos omnis sanguis iustus, qui effusus est super terram a sanguine Abel iusti usque ad sanguinem Zachariae filii Barachiae, quem occidistis inter templum et altare.
MATT|23|36|Amen dico vobis: Venient haec omnia super generationem istam.
MATT|23|37|Ierusalem, Ierusalem, quae occidis prophetas et lapidas eos, qui ad te missi sunt, quotiens volui congregare filios tuos, quemadmodum gallina congregat pullos suos sub alas, et noluistis!
MATT|23|38|Ecce relinquitur vobis domus vestra deserta!
MATT|23|39|Dico enim vobis: Non me videbitis amodo, donec dicatis: "Benedictus, qui venit in nomine Dominil" ".
MATT|24|1|Et egressus Iesus de templo ibat, et accesserunt discipuli eius, ut ostenderent ei aedificationes templi;
MATT|24|2|ipse autem respondens dixit eis: " Non videtis haec omnia? Amen dico vobis: Non relinquetur hic lapis super lapidem, qui non destruetur ".
MATT|24|3|Sedente autem eo super montem Oliveti, accesserunt ad eum discipuli secreto dicentes: " Dic nobis: Quando haec erunt, et quod signum adventus tui et consummationis saeculi? ".
MATT|24|4|Et respondens Iesus dixit eis: " Videte, ne quis vos seducat.
MATT|24|5|Multi enim venient in nomine meo dicentes: "Ego sum Christus", et multos seducent.
MATT|24|6|Audituri enim estis proelia et opiniones proeliorum. Videte, ne turbemini; oportet enim fieri, sed nondum est finis.
MATT|24|7|Consurget enim gens in gentem, et regnum in regnum, et erunt fames et terrae motus per loca;
MATT|24|8|haec autem omnia initia sunt dolorum.
MATT|24|9|Tunc tradent vos in tribulationem et occident vos, et eritis odio omnibus gentibus propter nomen meum.
MATT|24|10|Et tunc scandalizabuntur multi et invicem tradent et odio habebunt invicem;
MATT|24|11|et multi pseudoprophetae surgent et seducent multos.
MATT|24|12|Et, quoniam abundavit iniquitas, refrigescet caritas multorum;
MATT|24|13|qui autem permanserit usque in finem, hic salvus erit.
MATT|24|14|Et praedicabitur hoc evangelium regni in universo orbe in testimonium omnibus gentibus; et tunc veniet consummatio.
MATT|24|15|Cum ergo videritis abominationem desolationis, quae dicta est a Daniele propheta, stantem in loco sancto, qui legit, intellegat:
MATT|24|16|tunc qui in Iudaea sunt, fugiant ad montes;
MATT|24|17|qui in tecto, non descendat tollere aliquid de domo sua;
MATT|24|18|et, qui in agro, non revertatur tollere pallium suum.
MATT|24|19|Vae autem praegnantibus et nutrientibus in illis diebus!
MATT|24|20|Orate autem, ut non fiat fuga vestra hieme vel sabbato:
MATT|24|21|erit enim tunc tribulatio magna, qualis non fuit ab initio mundi usque modo neque fiet.
MATT|24|22|Et nisi breviati fuissent dies illi, non fieret salva omnis caro; sed propter electos breviabuntur dies illi.
MATT|24|23|Tunc si quis vobis dixerit: "Ecce hic Christus" aut: "Hic", nolite credere.
MATT|24|24|Surgent enim pseudochristi et pseudoprophetae et dabunt signa magna et prodigia, ita ut in errorem inducantur, si fieri potest, etiam electi.
MATT|24|25|Ecce praedixi vobis.
MATT|24|26|Si ergo dixerint vobis: "Ecce in deserto est", nolite exire; "Ecce in penetralibus", nolite credere;
MATT|24|27|sicut enim fulgur exit ab oriente et paret usque in occidentem, ita erit adventus Filii hominis.
MATT|24|28|Ubicumque fuerit corpus, illuc congregabuntur aquilae.
MATT|24|29|Statim autem post tribulationem dierum illorum, sol obscurabitur, et luna non dabit lumen suum, et stellae cadent de caelo, et virtutes caelorum commovebuntur.
MATT|24|30|Et tunc parebit signum Filii hominis in caelo, et tunc plangent omnes tribus terrae et videbunt Filium hominis venientem in nubibus caeli cum virtute et gloria multa;
MATT|24|31|et mittet angelos suos cum tuba magna, et congregabunt electos eius a quattuor ventis, a summis caelorum usque ad terminos eorum.
MATT|24|32|Ab arbore autem fici discite parabolam: cum iam ramus eius tener fuerit, et folia nata, scitis quia prope est aestas.
MATT|24|33|Ita et vos, cum videritis haec omnia, scitote quia prope est in ianuis.
MATT|24|34|Amen dico vobis: Non praeteribit haec generatio, donec omnia haec fiant.
MATT|24|35|Caelum et terra transibunt, verba vero mea non praeteribunt.
MATT|24|36|De die autem illa et hora nemo scit, neque angeli caelorum neque Filius, nisi Pater solus.
MATT|24|37|Sicut enim dies Noe, ita erit adventus Filii hominis.
MATT|24|38|Sicut enim erant in diebus ante diluvium comedentes et bibentes, nubentes et nuptum tradentes, usque ad eum diem, quo introivit in arcam Noe,
MATT|24|39|et non cognoverunt, donec venit diluvium et tulit omnes, ita erit et adventus Filii hominis.
MATT|24|40|Tunc duo erunt in agro: unus assumitur, et unus relinquitur;
MATT|24|41|duae molentes in mola: una assumitur, et una relinquitur.
MATT|24|42|Vigilate ergo, quia nescitis qua die Dominus vester venturus sit.
MATT|24|43|Illud autem scitote quoniam si sciret pater familias qua hora fur venturus esset, vigilaret utique et non sineret perfodi domum suam.
MATT|24|44|Ideo et vos estote parati, quia, qua nescitis hora, Filius hominis venturus est.
MATT|24|45|Quis putas est fidelis servus et prudens, quem constituit dominus supra familiam suam, ut det illis cibum in tempore?
MATT|24|46|Beatus ille servus, quem cum venerit dominus eius, invenerit sic facientem.
MATT|24|47|Amen dico vobis quoniam super omnia bona sua constituet eum.
MATT|24|48|Si autem dixerit malus servus ille in corde suo: "Moram facit dominus meus venire",
MATT|24|49|et coeperit percutere conservos suos, manducet autem et bibat cum ebriis,
MATT|24|50|veniet dominus servi illius in die, qua non sperat, et in hora, qua ignorat,
MATT|24|51|et dividet eum partemque eius ponet cum hypocritis; illic erit fletus et stridor dentium.
MATT|25|1|Tunc simile erit regnum cae lorum decem virginibus, quae accipientes lampades suas exierunt obviam sponso.
MATT|25|2|Quinque autem ex eis erant fatuae, et quinque prudentes.
MATT|25|3|Fatuae enim, acceptis lampadibus suis, non sumpserunt oleum secum;
MATT|25|4|prudentes vero acceperunt oleum in vasis cum lampadibus suis.
MATT|25|5|Moram autem faciente sponso, dormitaverunt omnes et dormierunt.
MATT|25|6|Media autem nocte clamor factus est: "Ecce sponsus! Exite obviam ei".
MATT|25|7|Tunc surrexerunt omnes virgines illae et ornaverunt lampades suas.
MATT|25|8|Fatuae autem sapientibus dixerunt: "Date nobis de oleo vestro, quia lampades nostrae exstinguuntur".
MATT|25|9|Responderunt prudentes dicentes: "Ne forte non sufficiat nobis et vobis, ite potius ad vendentes et emite vobis".
MATT|25|10|Dum autem irent emere, venit sponsus, et quae paratae erant, intraverunt cum eo ad nuptias; et clausa est ianua.
MATT|25|11|Novissime autem veniunt et reliquae virgines dicentes: "Domine, domine, aperi nobis".
MATT|25|12|At ille respondens ait: "Amen dico vobis: Nescio vos".
MATT|25|13|Vigilate itaque, quia nescitis diem neque horam.
MATT|25|14|Sicut enim homo peregre proficiscens vocavit servos suos et tradidit illis bona sua.
MATT|25|15|Et uni dedit quinque talenta, alii autem duo, alii vero unum, unicuique secundum propriam virtutem, et profectus est. Statim
MATT|25|16|abiit, qui quinque talenta acceperat, et operatus est in eis et lucratus est alia quinque;
MATT|25|17|similiter qui duo acceperat, lucratus est alia duo.
MATT|25|18|Qui autem unum acceperat, abiens fodit in terra et abscondit pecuniam domini sui.
MATT|25|19|Post multum vero temporis venit dominus servorum illorum et ponit rationem cum eis.
MATT|25|20|Et accedens, qui quinque talenta acceperat, obtulit alia quinque talenta dicens: "Domine, quinque talenta tradidisti mihi; ecce alia quinque superlucratus sum".
MATT|25|21|Ait illi dominus eius: "Euge, serve bone et fidelis. Super pauca fuisti fidelis; supra multa te constituam: intra in gaudium domini tui".
MATT|25|22|Accessit autem et qui duo talenta acceperat, et ait: "Domine, duo talenta tradidisti mihi; ecce alia duo lucratus sum".
MATT|25|23|Ait illi dominus eius: "Euge, serve bone et fidelis. Super pauca fuisti fidelis; supra multa te constituam: intra in gaudium domini tui".
MATT|25|24|Accedens autem et qui unum talentum acceperat, ait: "Domine, novi te quia homo durus es: metis, ubi non seminasti, et congregas, ubi non sparsisti;
MATT|25|25|et timens abii et abscondi talentum tuum in terra. Ecce habes, quod tuum est".
MATT|25|26|Respondens autem dominus eius dixit ei: "Serve male et piger! Sciebas quia meto, ubi non seminavi, et congrego, ubi non sparsi?
MATT|25|27|Oportuit ergo te mittere pecuniam meam nummulariis, et veniens ego recepissem, quod meum est cum usura.
MATT|25|28|Tollite itaque ab eo talentum et date ei, qui habet decem talenta:
MATT|25|29|omni enim habenti dabitur, et abundabit; ei autem, qui non habet, et quod habet, auferetur ab eo.
MATT|25|30|Et inutilem servum eicite in tenebras exteriores: illic erit fletus et stridor dentium".
MATT|25|31|Cum autem venerit Filius hominis in gloria sua, et omnes angeli cum eo, tunc sedebit super thronum gloriae suae.
MATT|25|32|Et congregabuntur ante eum omnes gentes; et separabit eos ab invicem, sicut pastor segregat oves ab haedis,
MATT|25|33|et statuet oves quidem a dextris suis, haedos autem a sinistris.
MATT|25|34|Tunc dicet Rex his, qui a dextris eius erunt: "Venite, benedicti Patris mei; possidete paratum vobis regnum a constitutione mundi.
MATT|25|35|Esurivi enim, et dedistis mihi manducare; sitivi, et dedistis mihi bibere; hospes eram, et collegistis me;
MATT|25|36|nudus, et operuistis me; infirmus, et visitastis me; in carcere eram, et venistis ad me".
MATT|25|37|Tunc respondebunt ei iusti dicentes: "Domine, quando te vidimus esurientem et pavimus, aut sitientem et dedimus tibi potum?
MATT|25|38|Quando autem te vidimus hospitem et collegimus, aut nudum et cooperuimus?
MATT|25|39|Quando autem te vidimus infirmum aut in carcere et venimus ad te?".
MATT|25|40|Et respondens Rex dicet illis: "Amen dico vobis: Quamdiu fecistis uni de his fratribus meis minimis, mihi fecistis".
MATT|25|41|Tunc dicet et his, qui a sinistris erunt: "Discedite a me, maledicti, in ignem aeternum, qui praeparatus est Diabolo et angelis eius.
MATT|25|42|Esurivi enim, et non dedistis mihi manducare; sitivi, et non dedistis mihi potum;
MATT|25|43|hospes eram, et non collegistis me; nudus, et non operuistis me; infirmus et in carcere, et non visitastis me".
MATT|25|44|Tunc respondebunt et ipsi dicentes: "Domine, quando te vidimus esurientem aut sitientem aut hospitem aut nudum aut infirmum vel in carcere et non ministravimus tibi?".
MATT|25|45|Tunc respondebit illis dicens: "Amen dico vobis: Quamdiu non fecistis uni de minimis his, nec mihi fecistis".
MATT|25|46|Et ibunt hi in supplicium aeternum, iusti autem in vitam aeternam ".
MATT|26|1|Et factum est, cum consum masset Iesus sermones hos omnes, dixit discipulis suis:
MATT|26|2|" Scitis quia post biduum Pascha fiet, et Filius hominis traditur, ut crucifigatur ".
MATT|26|3|Tunc congregati sunt principes sacerdotum et seniores populi in aulam principis sacerdotum, qui dicebatur Caiphas,
MATT|26|4|et consilium fecerunt, ut Iesum dolo tenerent et occiderent;
MATT|26|5|dicebant autem: " Non in die festo, ne tumultus fiat in populo ".
MATT|26|6|Cum autem esset Iesus in Bethania, in domo Simonis leprosi,
MATT|26|7|accessit ad eum mulier habens alabastrum unguenti pretiosi et effudit super caput ipsius recumbentis.
MATT|26|8|Videntes autem discipuli, indignati sunt dicentes: " Ut quid perditio haec?
MATT|26|9|Potuit enim istud venumdari multo et dari pauperibus ".
MATT|26|10|Sciens autem Iesus ait illis: " Quid molesti estis mulieri? Opus enim bonum operata est in me;
MATT|26|11|nam semper pauperes habetis vobiscum, me autem non semper habetis.
MATT|26|12|Mittens enim haec unguentum hoc supra corpus meum, ad sepeliendum me fecit.
MATT|26|13|Amen dico vobis: Ubicumque praedicatum fuerit hoc evangelium in toto mundo, dicetur et quod haec fecit in memoriam eius ".
MATT|26|14|Tunc abiit unus de Duodecim, qui dicebatur Iudas Iscariotes, ad principes sacerdotum
MATT|26|15|et ait: " Quid vultis mihi dare, et ego vobis eum tradam? ". At illi constituerunt ei triginta argenteos.
MATT|26|16|Et exinde quaerebat opportunitatem, ut eum traderet.
MATT|26|17|Prima autem Azymorum accesserunt discipuli ad Iesum dicentes: " Ubi vis paremus tibi comedere Pascha? ".
MATT|26|18|Ille autem dixit: " Ite in civitatem ad quendam et dicite ei: "Magister dicit: Tempus meum prope est; apud te facio Pascha cum discipulis meis" ".
MATT|26|19|Et fecerunt discipuli, sicut constituit illis Iesus, et paraverunt Pascha.
MATT|26|20|Vespere autem facto, discumbebat cum Duodecim.
MATT|26|21|Et edentibus illis, dixit: " Amen dico vobis: Unus vestrum me traditurus est ".
MATT|26|22|Et contristati valde, coeperunt singuli dicere ei: " Numquid ego sum, Domine? ".
MATT|26|23|At ipse respondens ait: " Qui intingit mecum manum in paropside, hic me tradet.
MATT|26|24|Filius quidem hominis vadit, sicut scriptum est de illo; vae autem homini illi, per quem Filius hominis traditur! Bonum erat ei, si natus non fuisset homo ille ".
MATT|26|25|Respondens autem Iudas, qui tradidit eum, dixit: " Numquid ego sum, Rabbi? ". Ait illi: " Tu dixisti ".
MATT|26|26|Cenantibus autem eis, accepit Iesus panem et benedixit ac fregit deditque discipulis et ait: " Accipite, comedite: hoc est corpus meum ".
MATT|26|27|Et accipiens calicem, gratias egit et dedit illis dicens: " Bibite ex hoc omnes:
MATT|26|28|hic est enim sanguis meus novi testamenti, qui pro multis effunditur in remissionem peccatorum.
MATT|26|29|Dico autem vobis: Non bibam amodo de hoc genimine vitis usque in diem illum, cum illud bibam vobiscum novum in regno Patris mei ".
MATT|26|30|Et hymno dicto, exierunt in montem Oliveti.
MATT|26|31|Tunc dicit illis Iesus: " Omnes vos scandalum patiemini in me in ista nocte. Scriptum est enim: "Percutiam pastorem, et dispergentur oves gregis".
MATT|26|32|Postquam autem resurrexero, praecedam vos in Galilaeam ".
MATT|26|33|Respondens autem Petrus ait illi: " Et si omnes scandalizati fuerint in te, ego numquam scandalizabor ".
MATT|26|34|Ait illi Iesus: " Amen dico tibi: In hac nocte, antequam gallus cantet, ter me negabis ".
MATT|26|35|Ait illi Petrus: " Etiam si oportuerit me mori tecum, non te negabo ". Similiter et omnes discipuli dixerunt.
MATT|26|36|Tunc venit Iesus cum illis in praedium, quod dicitur Gethsemani. Et dicit discipulis: " Sedete hic, donec vadam illuc et orem ".
MATT|26|37|Et assumpto Petro et duobus filiis Zebedaei, coepit contristari et maestus esse.
MATT|26|38|Tunc ait illis: " Tristis est anima mea usque ad mortem; sustinete hic et vigilate mecum ".
MATT|26|39|Et progressus pusillum, procidit in faciem suam orans et dicens: " Pater mi, si possibile est, transeat a me calix iste; verumtamen non sicut ego volo, sed sicut tu ".
MATT|26|40|Et venit ad discipulos et invenit eos dormientes; et dicit Petro: " Sic non potuistis una hora vigilare mecum?
MATT|26|41|Vigilate et orate, ut non intretis in tentationem; spiritus quidem promptus est, caro autem infirma ".
MATT|26|42|Iterum secundo abiit et oravit dicens: " Pater mi, si non potest hoc transire, nisi bibam illud, fiat voluntas tua ".
MATT|26|43|Et venit iterum et invenit eos dormientes: erant enim oculi eorum gravati.
MATT|26|44|Et relictis illis, iterum abiit et oravit tertio, eundem sermonem iterum dicens.
MATT|26|45|Tunc venit ad discipulos et dicit illis: " Dormite iam et requiescite; ecce appropinquavit hora, et Filius hominis traditur in manus peccatorum.
MATT|26|46|Surgite, eamus; ecce appropinquavit, qui me tradit ".
MATT|26|47|Et adhuc ipso loquente, ecce Iudas, unus de Duodecim, venit, et cum eo turba multa cum gladiis et fustibus, missi a principibus sacerdotum et senioribus populi.
MATT|26|48|Qui autem tradidit eum, dedit illis signum dicens: " Quemcumque osculatus fuero, ipse est; tenete eum! ".
MATT|26|49|Et confestim accedens ad Iesum dixit: " Ave, Rabbi! " et osculatus est eum.
MATT|26|50|Iesus autem dixit illi: " Amice, ad quod venisti! ". Tunc accesserunt et manus iniecerunt in Iesum et tenuerunt eum.
MATT|26|51|Et ecce unus ex his, qui erant cum Iesu, extendens manum exemit gladium suum et percutiens servum principis sacerdotum amputavit auriculam eius.
MATT|26|52|Tunc ait illi Iesus: " Converte gladium tuum in locum suum. Omnes enim, qui acceperint gladium, gladio peribunt.
MATT|26|53|An putas quia non possum rogare Patrem meum, et exhibebit mihi modo plus quam duodecim legiones angelorum?
MATT|26|54|Quomodo ergo implebuntur Scripturae quia sic oportet fieri? ".
MATT|26|55|In illa hora dixit Iesus turbis: " Tamquam ad latronem existis cum gladiis et fustibus comprehendere me? Cotidie sedebam docens in templo, et non me tenuistis ".
MATT|26|56|Hoc autem totum factum est, ut implerentur scripturae Prophetarum. Tunc discipuli omnes, relicto eo, fugerunt.
MATT|26|57|Illi autem tenentes Iesum duxerunt ad Caipham principem sacerdotum, ubi scribae et seniores convenerant.
MATT|26|58|Petrus autem sequebatur eum a longe usque in aulam principis sacerdotum; et ingressus intro sede bat cum ministris, ut videret finem.
MATT|26|59|Principes autem sacerdotum et omne concilium quaerebant falsum testimonium contra Iesum, ut eum morti traderent,
MATT|26|60|et non invenerunt, cum multi falsi testes accessissent. Novissime autem venientes duo
MATT|26|61|dixerunt: " Hic dixit: "Possum destruere templum Dei et post triduum aedificare illud" ".
MATT|26|62|Et surgens princeps sacerdotum ait illi: " Nihil respondes? Quid isti adversum te testificantur? ".
MATT|26|63|Iesus autem tacebat. Et princeps sacerdotum ait illi: " Adiuro te per Deum vivum, ut dicas nobis, si tu es Christus Filius Dei ".
MATT|26|64|Dicit illi Iesus: " Tu dixisti. Verumtamen dico vobis: Amodo videbitis Filium hominis sedentem a dextris Virtutis et venientem in nubibus caeli.
MATT|26|65|Tunc princeps sacerdotum scidit vestimenta sua dicens: " Blasphemavit! Quid adhuc egemus testibus? Ecce nunc audistis blasphemiam.
MATT|26|66|Quid vobis videtur? ". Illi autem respondentes dixerunt: " Reus est mortis! ".
MATT|26|67|Tunc exspuerunt in faciem eius et colaphis eum ceciderunt; alii autem palmas in faciem ei dederunt
MATT|26|68|dicentes: " Prophetiza nobis, Christe: Quis est, qui te percussit? ".
MATT|26|69|Petrus vero sedebat foris in atrio; et accessit ad eum una ancilla dicens: " Et tu cum Iesu Galilaeo eras! ".
MATT|26|70|At ille negavit coram omnibus dicens: " Nescio quid dicis! ".
MATT|26|71|Exeunte autem illo ad ianuam, vidit eum alia et ait his, qui erant ibi: Hic erat cum Iesu Nazareno! ".
MATT|26|72|Et iterum negavit cum iuramento: " Non novi hominem! ".
MATT|26|73|Post pusillum autem accesserunt, qui stabant, et dixerunt Petro: " Vere et tu ex illis es, nam et loquela tua manifestum te facit ".
MATT|26|74|Tunc coepit detestari et iurare: " Non novi hominem! ". Et continuo gallus cantavit;
MATT|26|75|et recordatus est Petrus verbi Iesu, quod dixerat: " Priusquam gallus cantet, ter me negabis ". Et egressus foras ploravit amare.
MATT|27|1|Mane autem facto, consi lium inierunt omnes princi pes sacerdotum et seniores populi adversus Iesum, ut eum morti traderent.
MATT|27|2|Et vinctum adduxerunt eum et tradiderunt Pilato praesidi.
MATT|27|3|Tunc videns Iudas, qui eum tradidit, quod damnatus esset, paenitentia ductus, rettulit triginta argenteos principibus sacerdotum et senioribus
MATT|27|4|dicens: " Peccavi tradens sanguinem innocentem ". At illi dixerunt: " Quid ad nos? Tu videris! ".
MATT|27|5|Et proiectis argenteis in templo, recessit et abiens laqueo se suspendit.
MATT|27|6|Principes autem sacerdotum, acceptis argenteis, dixerunt: " Non licet mittere eos in corbanam, quia pretium sanguinis est ".
MATT|27|7|Consilio autem inito, emerunt ex illis agrum Figuli in sepulturam peregrinorum.
MATT|27|8|Propter hoc vocatus est ager ille ager Sanguinis usque in hodiernum diem.
MATT|27|9|Tunc impletum est quod dictum est per Ieremiam prophetam di centem: " Et acceperunt triginta argenteos, pretium appretiati quem appretiaverunt a filiis Israel,
MATT|27|10|et dederunt eos in agrum Figuli, sicut constituit mihi Dominus ".
MATT|27|11|Iesus autem stetit ante praesidem; et interrogavit eum praeses dicens: Tu es Rex Iudaeorum? ". Dixit autem Iesus: " Tu dicis ".
MATT|27|12|Et cum accusaretur a principibus sacerdotum et senioribus, nihil respondit.
MATT|27|13|Tunc dicit illi Pilatus: " Non audis quanta adversum te dicant testimonia? ".
MATT|27|14|Et non respondit ei ad ullum verbum, ita ut miraretur praeses vehementer.
MATT|27|15|Per diem autem sollemnem consueverat praeses dimittere turbae unum vinctum, quem voluissent.
MATT|27|16|Habebant autem tunc vinctum insignem, qui dicebatur Barabbas.
MATT|27|17|Congregatis ergo illis dixit Pilatus: " Quem vultis dimittam vobis: Barabbam an Iesum, qui dicitur Christus? ".
MATT|27|18|Sciebat enim quod per invidiam tradidissent eum.
MATT|27|19|Sedente autem illo pro tribunali, misit ad illum uxor eius dicens: " Nihil tibi et iusto illi. Multa enim passa sum hodie per visum propter eum.
MATT|27|20|Principes autem sacerdotum et seniores persuaserunt turbis, ut peterent Barabbam, Iesum vero perderent.
MATT|27|21|Respondens autem praeses ait illis: " Quem vultis vobis de duobus dimittam? ". At illi dixerunt: " Barabbam! ".
MATT|27|22|Dicit illis Pilatus: " Quid igitur faciam de Iesu, qui dicitur Christus? ". Dicunt omnes: " Crucifigatur! ".
MATT|27|23|Ait autem: " Quid enim mali fecit? ". At illi magis clamabant dicentes: Crucifigatur! ".
MATT|27|24|Videns autem Pilatus quia nihil proficeret, sed magis tumultus fieret, accepta aqua, lavit manus coram turba dicens: " Innocens ego sum a sanguine hoc; vos videritis! ".
MATT|27|25|Et respondens universus populus dixit: " Sanguis eius super nos et super filios nostros ".
MATT|27|26|Tunc dimisit illis Barabbam; Iesum autem flagellatum tradidit, ut crucifigeretur.
MATT|27|27|Tunc milites praesidis suscipientes Iesum in praetorio congregaverunt ad eum universam cohortem.
MATT|27|28|Et exuentes eum, clamydem coccineam circumdederunt ei
MATT|27|29|et plectentes coronam de spinis posuerunt super caput eius et arundinem in dextera eius et, genu flexo ante eum, illudebant ei dicentes: " Ave, rex Iudaeorum! ".
MATT|27|30|Et exspuentes in eum acceperunt arundinem et percutiebant caput eius.
MATT|27|31|Et postquam illuserunt ei, exuerunt eum clamyde et induerunt eum vestimentis eius et duxerunt eum, ut crucifigerent.
MATT|27|32|Exeuntes autem invenerunt hominem Cyrenaeum nomine Simonem; hunc angariaverunt, ut tolleret crucem eius.
MATT|27|33|Et venerunt in locum, qui dicitur Golgotha, quod est Calvariae locus,
MATT|27|34|et dederunt ei vinum bibere cum felle mixtum; et cum gustasset, noluit bibere.
MATT|27|35|Postquam autem crucifixerunt eum, diviserunt vestimenta eius sortem mittentes
MATT|27|36|et sedentes servabant eum ibi.
MATT|27|37|Et imposuerunt super caput eius causam ipsius scriptam: " Hic est Iesus Rex Iudaeorum ".
MATT|27|38|Tunc crucifiguntur cum eo duo latrones: unus a dextris, et unus a sinistris.
MATT|27|39|Praetereuntes autem blasphemabant eum moventes capita sua
MATT|27|40|et dicentes: " Qui destruis templum et in triduo illud reaedificas, salva temetipsum; si Filius Dei es, descende de cruce! ".
MATT|27|41|Similiter et principes sacerdotum illudentes cum scribis et senioribus dicebant:
MATT|27|42|" Alios salvos fecit, seipsum non potest salvum facere. Rex Israel est; descendat nunc de cruce, et credemus in eum.
MATT|27|43|Confidit in Deo; liberet nunc, si vult eum. Dixit enim: "Dei Filius sum" ".
MATT|27|44|Idipsum autem et latrones, qui crucifixi erant cum eo, improperabant ei.
MATT|27|45|A sexta autem hora tenebrae factae sunt super universam terram usque ad horam nonam.
MATT|27|46|Et circa horam nonam clamavit Iesus voce magna dicens: " Eli, Eli, lema sabacthani? ", hoc est: " Deus meus, Deus meus, ut quid dereliquisti me?.
MATT|27|47|Quidam autem ex illic stantibus audientes dicebant: " Eliam vocat iste.
MATT|27|48|Et continuo currens unus ex eis acceptam spongiam implevit aceto et imposuit arundini et dabat ei bibere.
MATT|27|49|Ceteri vero dicebant: " Sine, videamus an veniat Elias liberans eum ".
MATT|27|50|Iesus autem iterum clamans voce magna emisit spiritum.
MATT|27|51|Et ecce velum templi scissum est a summo usque deorsum in duas partes, et terra mota est, et petrae scissae sunt;
MATT|27|52|et monumenta aperta sunt, et multa corpora sanctorum, qui dormierant, surrexerunt
MATT|27|53|et exeuntes de monumentis post resurrectionem eius venerunt in sanctam civitatem et apparuerunt multis.
MATT|27|54|Centurio autem et, qui cum eo erant custodientes Iesum, viso terrae motu et his, quae fiebant, timuerunt valde dicentes: " Vere Dei Filius erat iste! ".
MATT|27|55|Erant autem ibi mulieres multae a longe aspicientes, quae secutae erant Iesum a Galilaea ministrantes ei;
MATT|27|56|inter quas erat Maria Magdalene et Maria Iacobi et Ioseph mater et mater filiorum Zebedaei.
MATT|27|57|Cum sero autem factum esset, venit homo dives ab Arimathaea nomine Ioseph, qui et ipse discipulus erat Iesu.
MATT|27|58|Hic accessit ad Pilatum et petiit corpus Iesu. Tunc Pilatus iussit reddi.
MATT|27|59|Et accepto corpore, Ioseph involvit illud in sindone munda
MATT|27|60|et posuit illud in monumento suo novo, quod exciderat in petra, et advolvit saxum magnum ad ostium monumenti et abiit.
MATT|27|61|Erat autem ibi Maria Magdalene et altera Maria sedentes contra sepulcrum.
MATT|27|62|Altera autem die, quae est post Parascevem, convenerunt principes sacerdotum et pharisaei ad Pilatum
MATT|27|63|dicentes: " Domine, recordati sumus quia seductor ille dixit adhuc vivens: "Post tres dies resurgam".
MATT|27|64|Iube ergo custodiri sepulcrum usque in diem tertium, ne forte veniant discipuli eius et furentur eum et dicant plebi: "Surrexit a mortuis", et erit novissimus error peior priore ".
MATT|27|65|Ait illis Pilatus: " Habetis custodiam; ite, custodite, sicut scitis ".
MATT|27|66|Illi autem abeuntes munierunt sepulcrum, signantes lapidem, cum custodia.
MATT|28|1|Sero autem post sabbatum, cum illucesceret in primam sabbati, venit Maria Magdalene et altera Maria videre sepulcrum.
MATT|28|2|Et ecce terrae motus factus est magnus: angelus enim Domini descendit de caelo et accedens revolvit lapidem et sedebat super eum.
MATT|28|3|Erat autem aspectus eius sicut fulgur, et vestimentum eius candidum sicut nix.
MATT|28|4|Prae timore autem eius exterriti sunt custodes et facti sunt velut mortui.
MATT|28|5|Respondens autem angelus dixit mulieribus: " Nolite timere vos! Scio enim quod Iesum, qui crucifixus est, quaeritis.
MATT|28|6|Non est hic: surrexit enim, sicut dixit. Venite, videte locum, ubi positus erat.
MATT|28|7|Et cito euntes dicite discipulis eius: "Surrexit a mortuis et ecce praecedit vos in Galilaeam; ibi eum videbitis". Ecce dixi vobis ".
MATT|28|8|Et exeuntes cito de monumento cum timore et magno gaudio cucurrerunt nuntiare discipulis eius.
MATT|28|9|Et ecce Iesus occurrit illis dicens: " Avete ". Illae autem accesserunt et tenuerunt pedes eius et adoraverunt eum.
MATT|28|10|Tunc ait illis Iesus: " Nolite timere; ite, nuntiate fratribus meis, ut eant in Galilaeam et ibi me videbunt ".
MATT|28|11|Quae cum abiissent, ecce quidam de custodia venerunt in civitatem et nuntiaverunt principibus sacerdotum omnia, quae facta fuerant.
MATT|28|12|Et congregati cum senioribus, consilio accepto, pecuniam copiosam dederunt militibus
MATT|28|13|dicentes: " Dicite: "Discipuli eius nocte venerunt et furati sunt eum, nobis dormientibus".
MATT|28|14|Et si hoc auditum fuerit a praeside, nos suadebimus ei et securos vos faciemus ".
MATT|28|15|At illi, accepta pecunia, fecerunt, sicut erant docti. Et divulgatum est verbum istud apud Iudaeos usque in hodiernum diem.
MATT|28|16|Undecim autem discipuli abierunt in Galilaeam, in montem ubi constituerat illis Iesus,
MATT|28|17|et videntes eum adoraverunt; quidam autem dubitaverunt.
MATT|28|18|Et accedens Iesus locutus est eis dicens: " Data est mihi omnis potestas in caelo et in terra.
MATT|28|19|Euntes ergo docete omnes gentes, baptizantes eos in nomine Patris et Filii et Spiritus Sancti,
MATT|28|20|docentes eos servare omnia, quaecumque mandavi vobis. Et ecce ego vobiscum sum omnibus diebus usque ad consummationem saeculi ".
