1CHR|1|1|Адам, Сиф, Енос,
1CHR|1|2|Каинан, Малелеил, Иаред,
1CHR|1|3|Енох, Мафусал, Ламех,
1CHR|1|4|Ной, Сим, Хам и Иафет.
1CHR|1|5|Сыновья Иафета: Гомер, Магог, Мадай, Иаван, Фувал, Мешех и Фирас.
1CHR|1|6|Сыновья Гомера: Аскеназ, Рифат и Фогарма.
1CHR|1|7|Сыновья Иавана: Елиса, Фарсис, Киттим и Доданим.
1CHR|1|8|Сыновья Хама: Хуш, Мицраим, Фут и Ханаан.
1CHR|1|9|Сыновья Хуша: Сева, Хавила, Савта, Раама и Савтеха. Сыновья Раамы: Шева и Дедан.
1CHR|1|10|Хуш родил [также] Нимрода: сей начал быть сильным на земле.
1CHR|1|11|Мицраим родил: Лудима, Анамима, Легавима, Нафтухима,
1CHR|1|12|Патрусима, Каслухима, от которого произошли Филистимляне, и Кафторима.
1CHR|1|13|Ханаан родил Сидона, первенца своего, Хета,
1CHR|1|14|Иевусея, Аморрея, Гергесея,
1CHR|1|15|Евея, Аркея, Синея,
1CHR|1|16|Арвадея, Цемарея и Хамафея.
1CHR|1|17|Сыновья Сима: Елам, Ассур, Арфаксад, Луд, Арам, Уц, Хул, Гефер и Мешех.
1CHR|1|18|Арфаксад родил Салу, Сала же родил Евера.
1CHR|1|19|У Евера родились два сына: имя одному Фалек, потому что во дни его разделилась земля; имя брату его Иоктан.
1CHR|1|20|Иоктан родил Алмодада, Шалефа, Хацармавета, Иераха,
1CHR|1|21|Гадорама, Узала, Диклу,
1CHR|1|22|Евала, Авимаила, Шеву,
1CHR|1|23|Офира, Хавилу и Иовава. Все эти сыновья Иоктана.
1CHR|1|24|Сим, Арфаксад, Сала,
1CHR|1|25|Евер, Фалек, Рагав,
1CHR|1|26|Серух, Нахор, Фарра,
1CHR|1|27|Аврам, он же Авраам.
1CHR|1|28|Сыновья Авраама: Исаак и Измаил.
1CHR|1|29|Вот родословие их: первенец Измаилов Наваиоф, [за ним] Кедар, Адбеел, Мивсам,
1CHR|1|30|Мишма, Дума, Масса, Хадад, Фема,
1CHR|1|31|Иетур, Нафиш и Кедма. Это сыновья Измаиловы.
1CHR|1|32|Сыновья Хеттуры, наложницы Авраамовой: она родила Зимрана, Иокшана, Медана, Мадиана, Ишбака и Шуаха. Сыновья Иокшана: Шева и Дедан.
1CHR|1|33|Сыновья Мадиана: Ефа, Ефер, Ханох, Авида и Елдага. Все эти сыновья Хеттуры.
1CHR|1|34|И родил Авраам Исаака. Сыновья Исаака: Исав и Израиль.
1CHR|1|35|Сыновья Исава: Елифаз, Рагуил, Иеус, Иеглом и Корей.
1CHR|1|36|Сыновья Елифаза: Феман, Омар, Цефо, Гафам, Кеназ, Тимна, Амалика.
1CHR|1|37|Сыновья Рагуила: Нахаф, Зерах, Шамма и Миза.
1CHR|1|38|Сыновья Сеира: Лотан, Шовал, Цивеон, Ана, Дишон, Ецер и Дишан.
1CHR|1|39|Сыновья Лотана: Хори и Гемам; а сестра у Лотана: Фимна.
1CHR|1|40|Сыновья Шовала: Алеан, Манахаф, Евал, Шефо и Онам. Сыновья Цивеона: Аиа и Ана.
1CHR|1|41|Дети Аны: Дишон. Сыновья Дишона: Хемдан, Ешбан, Ифран и Херан.
1CHR|1|42|Сыновья Ецера: Билган, Зааван и Акан. Сыновья Дишана: Уц и Аран.
1CHR|1|43|Сии суть цари, царствовавшие в земле Едома, прежде нежели воцарился царь над сынами Израилевыми: Бела, сын Веора, и имя городу его – Дингава;
1CHR|1|44|и умер Бела, и воцарился по нем Иовав, сын Зераха, из Восоры.
1CHR|1|45|И умер Иовав, и воцарился по нем Хушам, из земли Феманитян.
1CHR|1|46|И умер Хушам, и воцарился по нем Гадад, сын Бедадов, который поразил Мадианитян на поле Моава; имя городу его: Авив.
1CHR|1|47|И умер Гадад, и воцарился по нем Самла, из Масреки.
1CHR|1|48|И умер Самла, и воцарился по нем Саул из Реховофа, [что] при реке.
1CHR|1|49|И умер Саул, и воцарился по нем Баал–Ханан, сын Ахбора.
1CHR|1|50|И умер Баал–Ханан, и воцарился по нем Гадар; имя городу его Пау; имя жене его Мегетавеель, дочь Матреда, дочь Мезагава.
1CHR|1|51|И умер Гадар. И были старейшины у Едома: старейшина Фимна, старейшина Алва, старейшина Иетеф,
1CHR|1|52|старейшина Оливема, старейшина Эла, старейшина Пинон,
1CHR|1|53|старейшина Кеназ, старейшина Феман, старейшина Мивцар,
1CHR|1|54|старейшина Магдиил, старейшина Ирам. Вот старейшины Идумейские.
1CHR|2|1|Вот сыновья Израиля: Рувим, Симеон, Левий, Иуда, Иссахар, Завулон,
1CHR|2|2|Дан, Иосиф, Вениамин, Неффалим, Гад и Асир.
1CHR|2|3|Сыновья Иуды: Ир, Онан и Силом, – трое родились у него от дочери Шуевой, Хананеянки. И был Ир, первенец Иудин, не благоугоден в очах Господа, и Он умертвил его.
1CHR|2|4|И Фамарь, невестка его, родила ему Фареса и Зару. Всех сыновей у Иуды было пятеро.
1CHR|2|5|Сыновья Фареса: Есром и Хамул.
1CHR|2|6|Сыновья Зары: Зимри, Ефан, Еман, Халкол и Дара; всех их пятеро.
1CHR|2|7|Сыновья Харми: Ахар, наведший беду на Израиля, нарушив заклятие.
1CHR|2|8|Сын Ефана: Азария.
1CHR|2|9|Сыновья Есрома, которые родились у него: Иерахмеил, Арам и Хелувай.
1CHR|2|10|Арам же родил Аминадава; Аминадав родил Наассона, князя сынов Иудиных;
1CHR|2|11|Наассон родил Салмона, Салмон родил Вооза;
1CHR|2|12|Вооз родил Овида, Овид родил Иессея;
1CHR|2|13|Иессей родил первенца своего Елиава, второго – Аминадава, третьего – Самму,
1CHR|2|14|четвертого – Нафанаила, пятого – Раддая,
1CHR|2|15|шестого – Оцема, седьмого – Давида.
1CHR|2|16|Сестры их: Саруия и Авигея. Сыновья Саруии: Авесса, Иоав и Азаил, трое.
1CHR|2|17|Авигея родила Амессу; отец же Амессы – Иефер, Измаильтянин.
1CHR|2|18|Халев, сын Есрома, родил от Азувы, жены [своей], и от Иериофы, и вот сыновья его: Иешер, Шовав и Ардон.
1CHR|2|19|И умерла Азува; и взял себе Халев Ефрафу, и она родила ему Хура.
1CHR|2|20|Хур родил Урия, Урий родил Веселиила.
1CHR|2|21|После Есром вошел к дочери Махира, отца Галаадова, и взял ее, будучи шестидесяти лет, и она родила ему Сегува.
1CHR|2|22|Сегув родил Иаира, и было у него двадцать три города в земле Галаадской.
1CHR|2|23|Но Гессуряне и Сирияне взяли у них селения Иаира, Кенаф и зависящие от него города, – шестьдесят городов. Все эти города сыновей Махира, отца Галаадова.
1CHR|2|24|По смерти Есрома в Халев–Ефрафе, жена Есромова, Авия, родила ему Ашхура, отца Фекои.
1CHR|2|25|Сыновья Иерахмеила, первенца Есромова, были: первенец Рам, [за] [ним] Вуна, Орен, Оцем и Ахия.
1CHR|2|26|Была у Иерахмеила и другая жена, имя ее Афара; она мать Онама.
1CHR|2|27|Сыновья Рама, первенца Иерахмеилова, были: Маац, Иамин и Екер.
1CHR|2|28|Сыновья Онама были: Шаммай и Иада. Сыновья Шаммая: Надав и Авишур.
1CHR|2|29|Имя жене Авишуровой Авихаиль, и она родила ему Ахбана и Молида.
1CHR|2|30|Сыновья Надава: Селед и Афаим. И умер Селед бездетным.
1CHR|2|31|Сын Афаима: Иший. Сын Ишия: Шешан. Сын Шешана: Ахлай.
1CHR|2|32|Сыновья Иады, брата Шаммаева: Иефер и Ионафан. Иефер умер бездетным.
1CHR|2|33|Сыновья Ионафана: Пелеф и Заза. Это сыновья Иерахмеила.
1CHR|2|34|У Шешана не было сыновей, а только дочери. У Шешана [был] раб, Египтянин, имя его Иарха;
1CHR|2|35|Шешан отдал дочь свою Иархе, рабу своему, в жену: и она родила ему Аттая.
1CHR|2|36|Аттай родил Нафана, Нафан родил Завада;
1CHR|2|37|Завад родил Ефлала, Ефлал родил Овида;
1CHR|2|38|Овид родил Иеуя, Иеуй родил Азарию;
1CHR|2|39|Азария родил Хелеца, Хелец родил Елеасу;
1CHR|2|40|Елеаса родил Сисмая, Сисмай родил Саллума;
1CHR|2|41|Саллум родил Иекамию, Иекамия родил Елишаму.
1CHR|2|42|Сыновья Халева, брата Иерахмеилова: Меша, первенец его, – он отец Зифа; и сыновья Мареши, отца Хеврона.
1CHR|2|43|Сыновья Хеврона: Корей и Таппуах, и Рекем и Шема.
1CHR|2|44|Шема родил Рахама, отца Иоркеамова, а Рекем родил Шаммая.
1CHR|2|45|Сын Шаммая Маон, а Маон – отец Беф–Цура.
1CHR|2|46|И Ефа, наложница Халевова, родила Харана, Моцу и Газеза. И Харан родил Газеза.
1CHR|2|47|Сыновья Иегдая: Регем, Иофам, Гешан, Пелет, Ефа и Шааф.
1CHR|2|48|Наложница Халевова, Мааха, родила Шевера и Фирхану;
1CHR|2|49|она же родила Шаафа, отца Мадманны, Шеву, отца Махбены и отца Гивеи. Дочь же Халева – Ахса.
1CHR|2|50|Вот сыновья Халева: сын Хур, первенец Ефрафы; Шовал, отец Кириаф–Иарима;
1CHR|2|51|Салма, отец Вифлеема; Хареф, отец Бефгадера.
1CHR|2|52|У Шовала, отца Кириаф–Иарима, были сыновья: Гарое, Хаци, Галменюхот.
1CHR|2|53|Племена Кириаф–Иарима: Ифрияне, Футияне, Шумафане и Мидраитяне. От сих произошли Цоряне и Ештаоляне.
1CHR|2|54|Сыновья Салмы: Вифлеемляне и Нетофафяне, венец дома Иоавова и половина Менухотян – Цоряне,
1CHR|2|55|и племена Соферийцев, живших в Иабеце, Тирейцы, Шимейцы, Сухайцы: это Кинеяне, происшедшие от Хамафа, отца Бетрехава.
1CHR|3|1|Сыновья Давида, родившиеся у него в Хевроне, были: первенец Амнон, от Ахиноамы Изреелитянки; второй – Далуия, от Авигеи Кармилитянки;
1CHR|3|2|третий – Авессалом, сын Маахи, дочери Фалмая, царя Гессурского; четвертый – Адония, сын Аггифы;
1CHR|3|3|пятый – Сафатия, от Авиталы; шестой – Ифреам, от Аглаи, жены его, –
1CHR|3|4|шесть родившихся у него в Хевроне; царствовал же он там семь лет и шесть месяцев; а тридцать три года царствовал в Иерусалиме.
1CHR|3|5|А сии родились у него в Иерусалиме: Шима, Шовав, Нафан и Соломон, четверо от Вирсавии, дочери Аммииловой;
1CHR|3|6|Ивхар, Елишама, Елифелет,
1CHR|3|7|Ногаг, Нефег, Иафиа,
1CHR|3|8|Елишама, Елиада и Елифелет – девятеро.
1CHR|3|9|[Вот] все сыновья Давида, кроме сыновей от наложниц. Сестра их Фамарь.
1CHR|3|10|Сын Соломона Ровоам; его сын Авия, его сын Аса, его сын Иосафат,
1CHR|3|11|его сын Иорам, его сын Охозия, его сын Иоас,
1CHR|3|12|его сын Амасия, его сын Азария, его сын Иофам,
1CHR|3|13|его сын Ахаз, его сын Езекия, его сын Манассия,
1CHR|3|14|его сын Амон, его сын Иосия.
1CHR|3|15|Сыновья Иосии: первенец Иоахаз, второй Иоаким, третий Седекия, четвертый Селлум.
1CHR|3|16|Сыновья Иоакима: Иехония, сын его; Седекия, сын его.
1CHR|3|17|Сыновья Иехонии: Асир, Салафиил, сын его;
1CHR|3|18|Малкирам, Федаия, Шенацар, Иезекия, Гошама и Савадия.
1CHR|3|19|И сыновья Федаии: Зоровавель и Шимей. Сыновья же Зоровавеля: Мешуллам и Ханания, и Шеломиф, сестра их,
1CHR|3|20|и еще пять: Хашува, Огел, Берехия, Хасадия и Иушав–Хесед.
1CHR|3|21|И сыновья Ханании: Фелатия и Исаия; его сын Рефаия, его сын Арнан, его сын Овадия, его сын Шехания.
1CHR|3|22|Сын Шехании: Шемаия; сыновья Шемаии: Хаттуш, Игеал, Бариах, Неария и Шафат, шестеро.
1CHR|3|23|Сыновья Неарии: Елиоенай, Езекия и Азрикам, трое.
1CHR|3|24|Сыновья Елиоеная: Годавьягу, Елеашив, Фелаия, Аккув, Иоханан, Делаия и Анани, семеро.
1CHR|4|1|Сыновья Иуды: Фарес, Есром, Харми, Хур и Шовал.
1CHR|4|2|Реаия, сын Шовала, родил Иахафа; Иахаф родил Ахума и Лагада: от них племена Цорян.
1CHR|4|3|И сии сыновья Етама: Изреель, Ишма и Идбаш, и сестра их, по имени Гацлелпони,
1CHR|4|4|Пенуел, отец Гедора, и Езер, отец Хуша. Вот сыновья Хура, первенца Ефрафы, отца Вифлеема.
1CHR|4|5|У Ахшура, отца Фекои, были две жены: Хела и Наара.
1CHR|4|6|И родила ему Наара Ахузама, Хефера, Фимни и Ахашфари; это сыновья Наары.
1CHR|4|7|Сыновья Хелы: Цереф, Цохар и Ефнан.
1CHR|4|8|Коц родил: Анува и Цовева и племена Ахархела, сына Гарумова.
1CHR|4|9|Иавис был знаменитее своих братьев. Мать дала ему имя Иавис, сказав: я родила его с болезнью.
1CHR|4|10|И воззвал Иавис к Богу Израилеву [и] сказал: о, если бы Ты благословил меня Твоим благословением, распространил пределы мои, и рука Твоя была со мною, охраняя [меня] от зла, чтобы я не горевал!.. И Бог ниспослал [ему], чего он просил.
1CHR|4|11|Хелув же, брат Шухи, родил Махира; он есть отец Ештона.
1CHR|4|12|Ештон родил Беф–Рафу, Пасеаха и Техинну, отца города Нааса; это жители Рехи.
1CHR|4|13|Сыновья Кеназа: Гофониил и Сераия. Сын Гофониила: Хафаф.
1CHR|4|14|Меонофай родил Офру, а Сераия родил Иоава, родоначальника долины плотников, потому что они были плотники.
1CHR|4|15|Сыновья Халева, сына Иефонниина: Ир, Ила и Наам. Сын Илы: Кеназ.
1CHR|4|16|Сыновья Иегаллелела: Зиф, Зифа, Фирия и Асареел.
1CHR|4|17|Сыновья Езры: Иефер, Меред, Ефер и Иалон; Иефер же родил Мерома, Шаммая и Ишбаха, отца Ешфемои.
1CHR|4|18|И жена его Иудия родила Иереда, отца Гедора, и Хевера, отца Сохо, и Иекуфиила, отца Занаоха. Это сыновья Бифьи, дочери фараоновой, которую взял Меред.
1CHR|4|19|Сыновья жены его Годии, сестры Нахама, отца Кеилы: Гарми и Ешфемоа – Маахатянин.
1CHR|4|20|Сыновья Симеона: Амнон, Ринна, Бенханан и Филон. Сыновья Ишия: Зохеф и Бензохеф.
1CHR|4|21|Сыновья Силома, сына Иудина: Ир, отец Лехи, и Лаеда, отец Мареши, и семейства выделывавших виссон, из дома Ашбеи,
1CHR|4|22|и Иоким, и жители Хозевы, и Иоаш и Сараф, которые имели владение в Моаве, и Иашувилехем; но это события древние.
1CHR|4|23|Они [были] горшечники, и жили при садах и в огородах; у царя для работ его жили они там.
1CHR|4|24|Сыновья Симеона: Немуил, Иамин, Иарив, Зерах и Саул.
1CHR|4|25|Шаллум сын его; его сын Мивсам; его сын Мишма.
1CHR|4|26|Сыновья Мишмы: Хаммуил, сын его; его сын Закур; его сын Шимей.
1CHR|4|27|У Шимея [было] шестнадцать сыновей и шесть дочерей; у братьев же его сыновей [было] немного, и все племя их не так было многочисленно, как племя сынов Иуды.
1CHR|4|28|Они жили в Вирсавии, Моладе, Хацаршуале,
1CHR|4|29|в Билге, в Ецеме, в Фоладе,
1CHR|4|30|в Вефуиле, в Хорме, в Циклаге,
1CHR|4|31|в Беф–Маркавофе, в Хацарсусиме, в Беф–Биреи и в Шаариме. Вот города их до царствования Давидова,
1CHR|4|32|с селами их: Етам, Аин, Риммон, Фокен и Ашан, – пять городов.
1CHR|4|33|И все селения их, которые находились вокруг сих городов до Ваала; вот места жительства их и родословия их.
1CHR|4|34|Мешовав, Иамлех и Иосия, сын Амассии,
1CHR|4|35|Иоил и Иегу, сын Иошиви, сына Сераии, сына Асиилова,
1CHR|4|36|Елиоенай, Иакова, Ишохаия, Асаия, Адиил, Ишимиил и Ванея,
1CHR|4|37|и Зиза, сын Шифия, сын Аллона, сын Иедаии, сын Шимрия, сын Шемаии.
1CHR|4|38|Сии поименованные [были] князьями племен своих, и дом отцов их разделился на многие отрасли.
1CHR|4|39|Они доходили до Герары и до восточной стороны долины, чтобы найти пастбища для стад своих;
1CHR|4|40|и нашли пастбища тучные и хорошие и землю обширную, спокойную и безопасную, потому что до них жило там [только] немного Хамитян.
1CHR|4|41|И пришли сии, по именам записанные, во дни Езекии, царя Иудейского, и перебили кочующих и оседлых, которые там находились, и истребили их навсегда и поселились на месте их, ибо там были пастбища для стад их.
1CHR|4|42|Из них же, из сынов Симеоновых, пошли к горе Сеир пятьсот человек: Фелатия, Неария, Рефаия и Узиил, сыновья Ишия, [были] во главе их;
1CHR|4|43|и побили уцелевший там остаток Амаликитян, и живут там до сего дня.
1CHR|5|1|Сыновья Рувима, первенца Израилева, – он первенец; но, когда осквернил он постель отца своего, первенство его отдано сыновьям Иосифа, сына Израилева, с тем однакож, чтобы не писаться им первородными;
1CHR|5|2|потому что Иуда был сильнейшим из братьев своих, и вождь от него, но первенство [перенесено] на Иосифа.
1CHR|5|3|Сыновья Рувима, первенца Израилева: Ханох, Фаллу, Хецрон и Харми.
1CHR|5|4|Сыновья Иоиля: Шемая, сын его; его сын Гог, его сын Шимей,
1CHR|5|5|его сын Миха, его сын Реаия, его сын Ваал,
1CHR|5|6|его сын Беера, которого отвел в плен Феглафелласар, царь Ассирийский. Он [был] князем Рувимлян.
1CHR|5|7|И братья его, по племенам их, по родословному списку их, были: главный Иеиель, потом Захария,
1CHR|5|8|и Бела, сын Азаза, сына Шемы, сына Иоиля. Он обитал в Ароере до Нево и Ваал–Меона;
1CHR|5|9|а к востоку он обитал до входа в пустыню, идущую от реки Евфрата, потому что стада их были многочисленны в земле Галаадской.
1CHR|5|10|Во дни Саула они вели войну с Агарянами, которые пали от рук их, а они стали жить в шатрах и по всей восточной стороне Галаада.
1CHR|5|11|Сыновья Гада жили напротив их в земле Васанской до Салхи:
1CHR|5|12|в Васане Иоиль был главный, Шафан второй, потом Иаанай и Шафат.
1CHR|5|13|Братьев их с семействами их было семь: Михаил, Мешуллам, Шева, Иорай, Иаакан, Зия и Евер.
1CHR|5|14|Вот сыновья Авихаила, сына Хурия, сына Иароаха, сына Галаада, сына Михаила, сына Иешишая, сына Иахдо, сына Буза.
1CHR|5|15|Ахи, сын Авдиила, сына Гуниева, [был] главою своего рода.
1CHR|5|16|Они жили в Галааде, в Васане и в зависящих от него городах и во всех окрестностях Сарона, до исхода их.
1CHR|5|17|Все они перечислены во дни Иоафама, царя Иудейского, и во дни Иеровоама, царя Израильского.
1CHR|5|18|У потомков Рувима и Гада и полуплемени Манассиина было людей воинственных, мужей носящих щит и меч, стреляющих из лука и приученных к битве, сорок четыре тысячи семьсот шестьдесят, выходящих на войну.
1CHR|5|19|И воевали они с Агарянами, Иетуром, Нафишем и Надавом.
1CHR|5|20|И подана была им помощь против них, и преданы были в руки их Агаряне и все, что у них было, потому что они во время сражения воззвали к Богу, и Он услышал их, за то, что они уповали на Него.
1CHR|5|21|И взяли они стада их: верблюдов пятьдесят тысяч, из мелкого скота двести пятьдесят тысяч, ослов две тысячи, и сто тысяч душ людей,
1CHR|5|22|потому что много пало убитых, так как от Бога было сражение сие. И жили они на месте их до переселения.
1CHR|5|23|Потомки полуколена Манассиина жили в той земле, от Васана до Ваал–Ермона и Сенира и до горы Ермона; и их было много.
1CHR|5|24|И вот главы поколений их: Ефер, Ишьи, Елиил, Азриил, Иеремия, Годавия и Иагдиил, мужи мощные, мужи именитые, главы родов своих.
1CHR|5|25|Но когда они согрешили против Бога отцов своих и стали блудно ходить вслед богов народов той земли, которых изгнал Бог от лица их,
1CHR|5|26|тогда Бог Израилев возбудил дух Фула, царя Ассирийского, и дух Феглафелласара, царя Ассирийского, и он выселил Рувимлян и Гадитян и половину колена Манассиина, и отвел их в Халах, и Хавор, и Ару, и на реку Гозан, – [где они] до сего дня.
1CHR|5|27|Сыновья Левия: Гирсон, Кааф и Мерари.
1CHR|5|28|Сыновья Каафа: Амрам, Ицгар, Хеврон и Узиил.
1CHR|5|29|Дети Амрама: Аарон, Моисей и Мариам. Сыновья Аарона: Надав, Авиуд, Елеазар и Ифамар.
1CHR|5|30|Елеазар родил Финееса, Финеес родил Авишуя;
1CHR|5|31|Авишуй родил Буккия, Буккий родил Озию;
1CHR|5|32|Озия родил Зерахию, Зерахия родил Мераиофа;
1CHR|5|33|Мераиоф родил Амарию, Амария родил Ахитува;
1CHR|5|34|Ахитув родил Садока, Садок родил Ахимааса;
1CHR|5|35|Ахимаас родил Азарию, Азария родил Иоанана;
1CHR|5|36|Иоанан родил Азарию, – это тот, который был священником в храме, построенном Соломоном в Иерусалиме.
1CHR|5|37|И родил Азария Амарию, Амария родил Ахитува;
1CHR|5|38|Ахитув родил Садока, Садок родил Селлума;
1CHR|5|39|Селлум родил Хелкию, Хелкия родил Азарию;
1CHR|5|40|Азария родил Сераию, Сераия родил Иоседека.
1CHR|5|41|Иоседек пошел [в плен], когда Господь переселил Иудеев и Иерусалимлян рукою Навуходоносора.
1CHR|6|1|Итак сыновья Левия: Гирсон, Кааф и Мерари.
1CHR|6|2|Вот имена сыновей Гирсоновых: Ливни и Шимей.
1CHR|6|3|Сыновья Каафа: Амрам, Ицгар, Хеврон и Узиил.
1CHR|6|4|Сыновья Мерари: Махли и Муши. Вот потомки Левия по родам их.
1CHR|6|5|У Гирсона: Ливни, сын его; Иахав, сын его; Зимма, сын его;
1CHR|6|6|Иоах, сын его; Иддо, сын его; Зерах, сын его; Иеафрай, сын его.
1CHR|6|7|Сыновья Каафа: Аминадав, сын его; Корей, сын его; Асир, сын его;
1CHR|6|8|Елкана, сын его; Евиасаф, сын его; Асир, сын его;
1CHR|6|9|Тахаф, сын его; Уриил, сын его; Узия, сын его; Саул, сын его.
1CHR|6|10|Сыновья Елканы: Амасай и Ахимоф.
1CHR|6|11|Елкана, сын его; Цофай, сын его; Нахаф, сын его;
1CHR|6|12|Елиаф, сын его; Иерохам, сын его, Елкана, сын его.
1CHR|6|13|Сыновья Самуила: первенец Иоиль, второй Авия.
1CHR|6|14|Сыновья Мерари: Махли; Ливни, сын его; Шимей, сын его; Уза, сын его;
1CHR|6|15|Шима, сын его; Хаггия, сын его; Асаия, сын его.
1CHR|6|16|Вот те, которых Давид поставил начальниками над певцами в доме Господнем, со времени поставления в нем ковчега.
1CHR|6|17|Они служили певцами пред скиниею собрания, доколе Соломон не построил дома Господня в Иерусалиме. И они становились на службу свою по уставу своему.
1CHR|6|18|Вот те, которые становились с сыновьями своими: из сыновей Каафовых – Еман певец, сын Иоиля, сын Самуила,
1CHR|6|19|сын Елканы, сын Иерохама, сын Елиила, сын Тоаха,
1CHR|6|20|сын Цуфа, сын Елканы, сын Махафа, сын Амасая,
1CHR|6|21|сын Елканы, сын Иоиля, сын Азарии, сын Цефании,
1CHR|6|22|сын Тахафа, сын Асира, сын Авиасафа, сын Корея,
1CHR|6|23|сын Ицгара, сын Каафа, сын Левия, сын Израиля;
1CHR|6|24|и брат его Асаф, стоявший на правой стороне его, – Асаф, сын Берехии, сын Шимы,
1CHR|6|25|сын Михаила, сын Ваасеи, сын Малхии,
1CHR|6|26|сын Ефния, сын Зераха, сын Адаии,
1CHR|6|27|сын Ефана, сын Зиммы, сын Шимия,
1CHR|6|28|сын Иахафа, сын Гирсона, сын Левия.
1CHR|6|29|А из сыновей Мерари, братьев их, – на левой стороне: Ефан, сын Кишия, сын Авдия, сын Маллуха,
1CHR|6|30|сын Хашавии, сын Амасии, сын Хелкии,
1CHR|6|31|сын Амция, сын Вания, сын Шемера,
1CHR|6|32|сын Махлия, сын Мушия, сын Мерари, сын Левия.
1CHR|6|33|Братья их левиты определены на всякие службы при доме Божием;
1CHR|6|34|Аарон же и сыновья его сожигали на жертвеннике всесожжения и на жертвеннике кадильном, и совершали всякое священнодействие во Святом Святых и для очищения Израиля во всем, как заповедал раб Божий Моисей.
1CHR|6|35|Вот сыновья Аарона: Елеазар, сын его; Финеес, сын его; Авиуд, сын его;
1CHR|6|36|Буккий, сын его; Уззий, сын его; Зерахия, сын его;
1CHR|6|37|Мераиоф, сын его; Амария, сын его; Ахитув, сын его;
1CHR|6|38|Садок, сын его; Ахимаас, сын его.
1CHR|6|39|И вот жилища их по селениям их в пределах их: сыновьям Аарона из племени Каафова, так как жребий выпал им,
1CHR|6|40|дали Хеврон, в земле Иудиной, и предместья его вокруг его;
1CHR|6|41|поля же сего города и села его отдали Халеву, сыну Иефонниину.
1CHR|6|42|Сыновьям Аарона дали также города убежищ: Хеврон и Ливну с их предместьями, Иаттир и Ештемоа и предместья его,
1CHR|6|43|и Хилен и предместья его, Давир и предместья его,
1CHR|6|44|и Ашан и предместья его, Вефсамис и предместья его,
1CHR|6|45|а от колена Вениаминова – Геву и предместья ее, и Аллемеф и предместья его, и Анафоф и предместья его: всех городов их в племенах их тринадцать городов.
1CHR|6|46|Остальным сыновьям Каафа, из семейств этого колена, [дано] по жребию десять городов из удела половины колена Манассиина.
1CHR|6|47|Сыновьям Гирсона по племенам их, от колена Иссахарова, и от колена Асирова, и от колена Неффалимова, и от колена Манассиина в Васане, [дано] тринадцать городов.
1CHR|6|48|Сыновьям Мерари по племенам их, от колена Рувимова, и от колена Гадова, и от колена Завулонова, [дано] по жребию двенадцать городов.
1CHR|6|49|Так дали сыны Израилевы левитам города и предместья их.
1CHR|6|50|Дали они по жребию от колена сыновей Иудиных, и от колена сыновей Симеоновых, и от колена сыновей Вениаминовых те города, которые они назвали по именам.
1CHR|6|51|Некоторым же племенам сыновей Каафовых даны были города от колена Ефремова.
1CHR|6|52|И дали им города убежищ: Сихем и предместья его на горе Ефремовой, и Гезер и предместья его,
1CHR|6|53|и Иокмеам и предместья его, и Беф–Орон и предместья его,
1CHR|6|54|и Аиалон и предместья его, и Гаф–Риммон и предместья его;
1CHR|6|55|от половины колена Манассиина – Анер и предместья его, Билеам и предместья его. Это поколению остальных сыновей Каафовых.
1CHR|6|56|Сыновьям Гирсона от племени полуколена Манассиина [дали] Голан в Васане и предместья его, и Аштароф и предместья его.
1CHR|6|57|От колена Иссахарова – Кедес и предместья его, Давраф и предместья его,
1CHR|6|58|и Рамоф и предместья его, и Анем и предместья его;
1CHR|6|59|от колена Асирова – Машал и предместья его, и Авдон и предместья его,
1CHR|6|60|и Хукок и предместья его, и Рехов и предместья его;
1CHR|6|61|от колена Неффалимова – Кедес в Галилее и предместья его, и Хаммон и предместья его, и Кириафаим и предместья его.
1CHR|6|62|А прочим сыновьям Мерариным – от колена Завулонова Риммон и предместья его, Фавор и предместья его.
1CHR|6|63|По ту сторону Иордана, против Иерихона, на восток от Иордана, от колена Рувимова [дали] Восор в пустыне и предместья его, и Иаацу и предместья ее,
1CHR|6|64|и Кедемоф и предместья его, и Мефааф и предместья его;
1CHR|6|65|от колена Гадова – Рамоф в Галааде и предместья его, и Маханаим и предместья его,
1CHR|6|66|и Есевон и предместья его, и Иазер и предместья его.
1CHR|7|1|Сыновья Иссахара: Фола, Фуа, Иашув и Шимрон, четверо.
1CHR|7|2|Сыновья Фолы: Уззий, Рефаия, Иериил, Иахмай, Ивсам и Самуил, главные в поколениях Фолы, люди воинственные в своих поколениях; число их во дни Давида было двадцать две тысячи и шестьсот.
1CHR|7|3|Сын Уззия: Израхия; а сыновья Израхии: Михаил, Овадиа, Иоиль и Ишшия, пятеро. Все они главные.
1CHR|7|4|У них, по родам их, по поколениям их, было готово к сражению войска тридцать шесть тысяч; потому что у них было много жен и сыновей.
1CHR|7|5|Братьев же их, во всех поколениях Иссахаровых, людей воинственных, было восемьдесят семь тысяч, внесенных в родословные записи.
1CHR|7|6|У Вениамина: Бела, Бехер и Иедиаил, трое.
1CHR|7|7|Сыновья Белы: Ецбон, Уззий, Уззиил, Иеримоф и Ири, пятеро, главы поколений, люди воинственные. В родословных списках записано их двадцать две тысячи тридцать четыре.
1CHR|7|8|Сыновья Бехера: Земира, Иоаш, Елиезер, Елиоенай, Омри, Иремоф, Авия, Анафоф и Алемеф: все эти сыновья Бехера.
1CHR|7|9|В родословных списках записано их по родам их, по главам поколений, людей воинственных – двадцать тысяч и двести.
1CHR|7|10|Сын Иедиаила: Билган. Сыновья Билгана: Иеус, Вениамин, Егуд, Хенаана, Зефан, Фарсис и Ахишахар.
1CHR|7|11|Все эти сыновья Иедиаила были главами поколений, люди воинственные; семнадцать тысяч и двести было выходящих на войну.
1CHR|7|12|И Шупим и Хупим, сыновья Ира; Хушим, сын Ахера;
1CHR|7|13|сыновья Неффалима: Иахцеил, Гуни, Иецер и Шиллем, дети Валлы.
1CHR|7|14|Сыновья Манассии: Асриил, которого родила наложница его Арамеянка; она же родила Махира, отца Галаадова.
1CHR|7|15|Махир взял в жену сестру Хупима и Шупима, – имя сестры их Мааха; имя второму Салпаад. У Салпаада были [только] дочери.
1CHR|7|16|Мааха, жена Махирова, родила сына и нарекла ему имя Кереш, а имя брату его Шереш. Сыновья его: Улам и Рекем.
1CHR|7|17|Сын Улама: Бедан. Вот сыновья Галаада, сына Махира, сына Манассиина.
1CHR|7|18|Сестра его Молехеф родила Ишгода, Авиезера и Махлу.
1CHR|7|19|Сыновья Шемиды были: Ахиан, Шехем, Ликхи и Аниам.
1CHR|7|20|Сыновья Ефрема: Шутелах, и Беред, сын его, и Фахаф, сын его, и Елеада, сын его, и Фахаф, сын его,
1CHR|7|21|и Завад, сын его, и Шутелах, сын его, и Езер и Елеад. И убили их жители Гефа, уроженцы той земли, за то, что они пошли захватить стада их.
1CHR|7|22|И плакал о них Ефрем, отец их, много дней, и приходили братья его утешать его.
1CHR|7|23|Потом он вошел к жене своей, и она зачала и родила сына, и он нарек ему имя: Берия, потому что несчастье постигло дом его.
1CHR|7|24|И дочь у него [была] Шеера. Она построила Беф–Орон нижний и верхний и Уззен–Шееру.
1CHR|7|25|И Рефай, сын его, и Решеф, и Фелах, сын его, и Фахан, сын его,
1CHR|7|26|Лаедан, сын его, Аммиуд, сын его, Елишама, сын его,
1CHR|7|27|Нон, сын его, Иисус, сын его.
1CHR|7|28|Владения их и места жительства их [были]: Вефиль и зависящие от него города; к востоку Нааран, к западу Гезер и зависящие от него города; Сихем и зависящие от него города до Газы и зависящих от нее городов.
1CHR|7|29|А со стороны сыновей Манассииных: Беф–Сан и зависящие от него города, Фаанах и зависящие от него города, Мегиддо и зависящие от него города, Дор и зависящие от него города. В них жили сыновья Иосифа, сына Израилева.
1CHR|7|30|Сыновья Асира: Имна, Ишва, Ишви и Берия, и сестра их Серах.
1CHR|7|31|Сыновья Берии: Хевер и Малхиил. Он отец Бирзаифа.
1CHR|7|32|Хевер родил Иафлета, Шомера и Хофама, и Шую, сестру их.
1CHR|7|33|Сыновья Иафлета: Пасах, Бимгал и Ашваф. Вот сыновья Иафлета.
1CHR|7|34|Сыновья Шемера: Ахи, Рохга, Ихубба и Арам.
1CHR|7|35|Сыновья Гелема, брата его: Цофах, Имна, Шелеш и Амал.
1CHR|7|36|Сыновья Цофаха: Суах, Харнефер, Шуал, Бери, Имра,
1CHR|7|37|Бецер, Год, Шамма, Шилша, Ифран и Беера.
1CHR|7|38|Сыновья Иефера: Иефунни, Фиспа и Ара.
1CHR|7|39|Сыновья Уллы: Арах, Ханниил и Риция.
1CHR|7|40|Все эти сыновья Асира, главы поколений, люди отборные, воинственные, главные начальники. Записано у них в родословных списках в войске, для войны, по счету двадцать шесть тысяч человек.
1CHR|8|1|Вениамин родил Белу, первенца своего, второго Ашбела, третьего Ахрая,
1CHR|8|2|четвертого Ноху и пятого Рафу.
1CHR|8|3|Сыновья Белы были: Аддар, Гера, Авиуд,
1CHR|8|4|Авишуа, Нааман, Ахоах,
1CHR|8|5|Гера, Шефуфан и Хурам.
1CHR|8|6|И вот сыновья Егуда, которые были главами родов, живших в Геве и переселенных в Манахаф:
1CHR|8|7|Нааман, Ахия и Гера, который переселил их; он родил Уззу и Ахихуда.
1CHR|8|8|Шегараим родил детей в земле Моавитской после того, как отпустил от [себя] Хушиму и Баару, жен своих.
1CHR|8|9|И родил он от Ходеши, жены своей, Иовава, Цивию, Мешу, Малхама,
1CHR|8|10|Иеуца, Шахию и Мирму: вот сыновья его, главы поколений.
1CHR|8|11|От Хушимы родил он Авитува и Елпаала.
1CHR|8|12|Сыновья Елпаала: Евер, Мишам и Шемер, который построил Оно и Лод и зависящие от него города, –
1CHR|8|13|и Берия и Шема. Они были главами поколений жителей Аиалона. Они выгнали жителей Гефа.
1CHR|8|14|Ахио, Шашак, Иремоф,
1CHR|8|15|Зевадия, Арад, Едер,
1CHR|8|16|Михаил, Ишфа и Иоха – сыновья Берии.
1CHR|8|17|Зевадия, Мешуллам, Хизкий, Хевер,
1CHR|8|18|Ишмерай, Излия и Иовав – сыновья Елпаала.
1CHR|8|19|Иаким, Зихрий, Завдий,
1CHR|8|20|Елиенай, Цилфай, Елиил,
1CHR|8|21|Адаия, Бераия и Шимраф – сыновья Шимея.
1CHR|8|22|Ишпан, Евер, Елиил,
1CHR|8|23|Авдон, Зихрий, Ханан,
1CHR|8|24|Ханания, Елам, Антофия,
1CHR|8|25|Ифдия и Фенуил – сыновья Шашака.
1CHR|8|26|Шамшерай, Шехария, Афалия,
1CHR|8|27|Иаарешия, Елия и Зихрий, сыновья Иерохама.
1CHR|8|28|Это главы поколений, в родах своих главные. Они жили в Иерусалиме.
1CHR|8|29|В Гаваоне жили: отец Гаваонитян, – имя жены его Мааха, –
1CHR|8|30|и сын его, первенец Авдон, [за ним] Цур, Кис, Ваал, Надав,
1CHR|8|31|Гедор, Ахио, Зехер и Миклоф.
1CHR|8|32|Миклоф родил Шимея. И они подле братьев своих жили в Иерусалиме, вместе с братьями своими.
1CHR|8|33|Нер родил Киса; Кис родил Саула; Саул родил Иоанафана, Мелхисуя, Авинадава и Ешбаала.
1CHR|8|34|Сын Ионафана Мериббаал; Мериббаал родил Миху.
1CHR|8|35|Сыновья Михи: Пифон, Мелег, Фаарея и Ахаз.
1CHR|8|36|Ахаз родил Иоиадду; Иоиадда родил Алемефа, Азмавефа и Замврия; Замврий родил Моцу;
1CHR|8|37|Моца родил Бинею. Рефаия, сын его; Елеаса, сын его; Ацел, сын его.
1CHR|8|38|У Ацела шесть сыновей, и вот имена их: Азрикам, Бохру, Исмаил, Шеария, Овадия и Ханан; все они сыновья Ацела.
1CHR|8|39|Сыновья Ешека, брата его: Улам, первенец его, второй Иеуш, третий Елифелет.
1CHR|8|40|Сыновья Улама были люди воинственные, стрелявшие из лука, имевшие много сыновей и внуков: сто пятьдесят. Все они от сынов Вениамина.
1CHR|9|1|Так были перечислены по родам своим все Израильтяне, и вот они записаны в книге царей Израильских. Иудеи же за беззакония свои переселены в Вавилон.
1CHR|9|2|Первые жители, которые [жили] во владениях своих, по городам Израильским, были Израильтяне, священники, левиты и нефинеи.
1CHR|9|3|В Иерусалиме жили некоторые из сынов Иудиных и из сынов Вениаминовых, и из сынов Ефремовых и Манассииных:
1CHR|9|4|Уфай, сын Аммиуда, сын Омри, сын Имрия, сын Вания, – из сыновей Фареса, сына Иудина;
1CHR|9|5|из сыновей Шилона – Асаия первенец и сыновья его;
1CHR|9|6|из сыновей Зары – Иеуил и братья их, – шестьсот девяносто;
1CHR|9|7|из сыновей Вениаминовых Саллу, сын Мешуллама, сын Годавии, сын Гассенуи;
1CHR|9|8|и Ивния, сын Иерохама, и Эла, сын Уззия, сына Михриева, и Мешуллам, сын Шефатии, сына Регуила, сына Ивнии,
1CHR|9|9|и братья их, по родам их: девятьсот пятьдесят шесть, – все сии мужи были главы родов в поколениях своих.
1CHR|9|10|А из священников: Иедаия, Иоиарив, Иахин,
1CHR|9|11|и Азария, сын Хелкии, сын Мешуллама, сын Садока, сын Мераиофа, сын Ахитува, начальствующий в доме Божием;
1CHR|9|12|и Адаия, сын Иерохама, сын Пашхура, сын Малхии; и Маасай, сын Адиела, сын Иахзера, сын Мешуллама, сын Мешиллемифа, сын Иммера;
1CHR|9|13|и братья их, главы родов своих: тысяча семьсот шестьдесят, – люди отличные в деле служения в доме Божием.
1CHR|9|14|А из левитов: Шемаия, сын Хашува, сын Азрикама, сын Хашавии, – из сыновей Мерариных;
1CHR|9|15|и Вакбакар, Хереш, Галал, и Матфания, сын Михи, сын Зихрия, сын Асафа;
1CHR|9|16|и Овадия, сын Шемаии, сын Галала, сын Идифуна, и Берехия, сын Асы, сын Елканы, живший в селениях Нетофафских.
1CHR|9|17|А привратники: Шаллум, Аккуб, Талмон и Ахиман, и братья их; Шаллум [был] главным.
1CHR|9|18|И доныне сии привратники у ворот царских, к востоку, содержат стражу сынов Левииных.
1CHR|9|19|Шаллум, сын Коре, сын Евиасафа, сын Корея, и братья его из рода его, Кореяне, по делу служения своего, были стражами у порогов скинии, а отцы их охраняли вход в стан Господень.
1CHR|9|20|Финеес, сын Елеазаров, был прежде начальником над ними, и Господь был с ним.
1CHR|9|21|Захария, сын Мешелемии, [был] привратником у дверей скинии собрания.
1CHR|9|22|Всех их, выбранных в привратники к порогам, было двести двенадцать. Они внесены в список по селениям своим. Их поставил Давид и Самуил–прозорливец за верность их.
1CHR|9|23|И они и сыновья их были на страже у ворот дома Господня, при доме скинии.
1CHR|9|24|На четырех сторонах находились привратники: на восточной, западной, северной и южной.
1CHR|9|25|Братья же их жили в селениях своих, приходя к ним от времени до времени на семь дней.
1CHR|9|26|Сии четыре начальника привратников, левиты, были в доверенности; они же были приставлены к жилищам и к сокровищам дома Божия.
1CHR|9|27|Вокруг дома Божия они и ночь проводили, потому что на них [лежало] охранение, и они должны были каждое утро отпирать двери.
1CHR|9|28|[Одни] из них были приставлены к служебным сосудам, так что счетом принимали их и счетом выдавали.
1CHR|9|29|[Другим] из них поручена была прочая утварь и все священные потребности: мука лучшая, и вино, и елей, и ладан, и благовония.
1CHR|9|30|А из сыновей священнических [некоторые] составляли миро из веществ благовонных.
1CHR|9|31|Маттафии из левитов, – он первенец Селлума Кореянина, – вверено было приготовляемое на сковородах.
1CHR|9|32|[Некоторым] из братьев их, из сынов Каафовых, поручено было [заготовление] хлебов предложения, чтобы представлять [их] каждую субботу.
1CHR|9|33|Певцы же, главные в поколениях левитских, в комнатах храма свободны были от занятий, потому что день и ночь они обязаны были [заниматься] искусством [своим].
1CHR|9|34|Это главы поколений левитских, в родах своих главные. Они жили в Иерусалиме.
1CHR|9|35|В Гаваоне жили: отец Гаваонитян Иеил, – имя жены его Мааха,
1CHR|9|36|и сын его первенец Авдон, [за ним] Цур, Кис, Ваал, Нер, Надав,
1CHR|9|37|Гедор, Ахио, Захария и Миклоф.
1CHR|9|38|Миклоф родил Шимеама. И они подле братьев своих жили в Иерусалиме вместе с братьями своими.
1CHR|9|39|Нер родил Киса, Кис родил Саула, Саул родил Ионафана, Мелхисуя, Авинадава и Ешбаала.
1CHR|9|40|Сын Ионафана Мериббаал; Мериббаал родил Миху.
1CHR|9|41|Сыновья Михи: Пифон, Мелех, Фарей [и Ахаз].
1CHR|9|42|Ахаз родил Иаеру; Иаера родил Алемефа, Азмавефа и Замврия; Замврий родил Моцу;
1CHR|9|43|Моца родил Бинею: Рефаия, сын его; Елеаса, сын его; Ацел, сын его.
1CHR|9|44|У Ацела шесть сыновей, и вот имена их: Азрикам, Бохру, Исмаил, Шеария, Овадия и Ханан. Это сыновья Ацела.
1CHR|10|1|Филистимляне воевали с Израилем, и побежали Израильтяне от Филистимлян, и падали пораженные на горе Гелвуе.
1CHR|10|2|И погнались Филистимляне за Саулом и сыновьями его, и убили Филистимляне Ионафана и Авинадава и Мелхисуя, сыновей Сауловых.
1CHR|10|3|Сражение против Саула усилилось, и стрелки устремились на него, так что он изранен был стрелками.
1CHR|10|4|И сказал Саул оруженосцу своему: обнажи меч твой и заколи меня им, чтобы не пришли эти необрезанные и не надругались надо мною. Но оруженосец не решился, потому что очень испугался. Тогда Саул взял меч и пал на него.
1CHR|10|5|Оруженосец его, увидев, что Саул умер, и сам пал на меч и умер.
1CHR|10|6|И умер Саул, и три сына его, и весь дом его вместе с ним умер.
1CHR|10|7|Когда увидели Израильтяне, которые были в долине, что все бегут и что Саул и сыновья его умерли, то оставили города свои и разбежались; а Филистимляне пришли и поселились в них.
1CHR|10|8|На другой день пришли Филистимляне обирать убитых, и нашли Саула и сыновей его, павших на горе Гелвуйской,
1CHR|10|9|и раздели его, и сняли с него голову его и оружие его, и послали по земле Филистимской, чтобы возвестить [о сем] пред идолами их и пред народом.
1CHR|10|10|И положили оружие его в капище богов своих, и голову его воткнули в доме Дагона.
1CHR|10|11|И услышал весь Иавис Галаадский все, что сделали Филистимляне с Саулом.
1CHR|10|12|И поднялись все люди сильные, взяли тело Саулово и тела сыновей его, и принесли их в Иавис, и похоронили кости их под дубом в Иависе, и постились семь дней.
1CHR|10|13|Так умер Саул за свое беззаконие, которое он сделал пред Господом, за то, что не соблюл слова Господня и обратился к волшебнице с вопросом,
1CHR|10|14|а не взыскал Господа. [За то] Он и умертвил его, и передал царство Давиду, сыну Иессееву.
1CHR|11|1|И собрались все Израильтяне к Давиду в Хеврон и сказали: вот, мы кость твоя и плоть твоя;
1CHR|11|2|и вчера, и третьего дня, когда еще Саул был царем, ты выводил и вводил Израиля, и Господь Бог твой сказал тебе: "ты будешь пасти народ Мой, Израиля и ты будешь вождем народа Моего Израиля".
1CHR|11|3|И пришли все старейшины Израилевы к царю в Хеврон, и заключил с ними Давид завет в Хевроне пред лицем Господним; и они помазали Давида в царя над Израилем, по слову Господню, чрез Самуила.
1CHR|11|4|И пошел Давид и весь Израиль к Иерусалиму, то есть к Иевусу. А там были Иевусеи, жители той земли.
1CHR|11|5|И сказали жители Иевуса Давиду: не войдешь сюда. Но Давид взял крепость Сион; это город Давидов.
1CHR|11|6|И сказал Давид: кто прежде всех поразит Иевусеев, тот будет главою и военачальником. И взошел прежде всех Иоав, сын Саруи, и сделался главою.
1CHR|11|7|Давид жил в той крепости, потому и называли ее городом Давидовым.
1CHR|11|8|И он обстроил город кругом, [начиная] от Милло, всю окружность, а Иоав возобновил остальные [части] города.
1CHR|11|9|И преуспевал Давид, и возвышался более и более, и Господь Саваоф [был] с ним.
1CHR|11|10|Вот главные из сильных у Давида, которые крепко подвизались с ним в царстве его, вместе со всем Израилем, чтобы воцарить его, по слову Господню, над Израилем,
1CHR|11|11|и вот число храбрых, которые были у Давида: Иесваал, сын Ахамани, главный из тридцати. Он поднял копье свое на триста человек и поразил их в один раз.
1CHR|11|12|По нем Елеазар, сын Додо Ахохиянина, из трех храбрых:
1CHR|11|13|он был с Давидом в Фасдамиме, куда Филистимляне собрались на войну. Там часть поля была засеяна ячменем, и народ побежал от Филистимлян;
1CHR|11|14|но они стали среди поля, сберегли его и поразили Филистимлян. И даровал Господь спасение великое!
1CHR|11|15|Трое сих главных из тридцати вождей взошли на скалу к Давиду, в пещеру Одоллам, когда стан Филистимлян был расположен в долине Рефаимов.
1CHR|11|16|Давид тогда был в укрепленном месте, а охранное войско Филистимлян было тогда в Вифлееме.
1CHR|11|17|И сильно захотелось [пить] Давиду, и он сказал: кто напоит меня водою из колодезя Вифлеемского, что у ворот?
1CHR|11|18|Тогда эти трое пробились сквозь стан Филистимский и почерпнули воды из колодезя Вифлеемского, что у ворот, и взяли, и принесли Давиду. Но Давид не захотел пить ее и вылил ее во славу Господа,
1CHR|11|19|и сказал: сохрани меня Господь, чтоб я сделал это! Стану ли я пить кровь мужей сих, полагавших души свои! Ибо с опасностью собственной жизни они принесли [воду]. И не захотел пить ее. Вот что сделали трое этих храбрых.
1CHR|11|20|И Авесса, брат Иоава, был главным из трех: он убил копьем своим триста человек, и был в славе у тех троих.
1CHR|11|21|Из трех он был знатнейшим и был начальником; но с теми тремя не равнялся.
1CHR|11|22|Ванея, сын Иодая, мужа храброго, великий по делам, из Кавцеила: он поразил двух Ариилов Моавитских; он же сошел и убил льва во рве, в снежное время;
1CHR|11|23|он же убил Египтянина, человека ростом в пять локтей: в руке Египтянина было копье, как навой у ткачей, а он подошел к нему с палкою и, вырвав копье из руки Египтянина, убил его его же копьем:
1CHR|11|24|вот что сделал Ванея, сын Иодая. И он был в славе у тех троих храбрых;
1CHR|11|25|он был знатнее тридцати, но с тремя не равнялся, и Давид поставил его ближайшим исполнителем своих приказаний.
1CHR|11|26|А главные из воинов: Асаил, брат Иоава; Елханан, сын Додо, из Вифлеема;
1CHR|11|27|Шамма Гародитянин; Херец Пелонитянин;
1CHR|11|28|Ира, сын Икеша, Фекоитянин; Евиезер Анафофянин;
1CHR|11|29|Сивхай Хушатянин; Илай Ахохиянин;
1CHR|11|30|Магарай Нетофафянин; Хелед, сын Вааны, Нетофафянин;
1CHR|11|31|Иттай, сын Рибая, из Гивы Вениаминовой; Ванея Пирафонянин;
1CHR|11|32|Хурай из Нагале–Гааша; Авиел из Аравы;
1CHR|11|33|Азмавеф Бахарумиянин; Елияхба Шаалбонянин.
1CHR|11|34|Сыновья Гашема Гизонитянина: Ионафан, сын Шаге, Гараритянин;
1CHR|11|35|Ахиам, сын Сахара, Гараритянин; Елифал, сын Уры;
1CHR|11|36|Хефер из Махеры; Ахиа Пелонитянин;
1CHR|11|37|Хецрой Кармилитянин; Наарай, сын Езбая;
1CHR|11|38|Иоиль, брат Нафана; Мивхар, сын Гагрия;
1CHR|11|39|Целек Аммонитянин; Нахарай Берофянин, оруженосец Иоава, сына Саруи;
1CHR|11|40|Ира Ифриянин; Гареб Ифриянин;
1CHR|11|41|Урия Хеттеянин; Завад, сын Ахлая;
1CHR|11|42|Адина, сын Шизы, Рувимлянин, глава Рувимлян, и у него [было] тридцать;
1CHR|11|43|Ханан, сын Маахи; Иосафат Мифниянин;
1CHR|11|44|Уззия Аштерофянин; Шама и Иеиел, сыновья Хофама Ароерянина;
1CHR|11|45|Иедиаел, сын Шимрия, и Иоха, брат его, Фициянин;
1CHR|11|46|Елиел из Махавима, и Иеривай и Иошавия, сыновья Елнаама, и Ифма Моавитянин;
1CHR|11|47|Елиел, Овед и Иасиел из Мецоваи.
1CHR|12|1|И сии также пришли к Давиду в Секелаг, когда он еще укрывался от Саула, сына Кисова, и были из храбрых, помогавших в сражении.
1CHR|12|2|Вооруженные луком, правою и левою рукою [бросавшие] каменья и [стрелявшие] стрелами из лука, – из братьев Саула, от Вениамина:
1CHR|12|3|главный Ахиезер, за ним Иоас, сыновья Шемаи, из Гивы; Иезиел и Фелет, сыновья Азмавефа; Бераха и Иегу из Анафофа;
1CHR|12|4|Ишмаия Гаваонитянин, храбрый из тридцати и [начальствовавший] над тридцатью;
1CHR|12|5|Иеремия, Иахазиил, Иоханан и Иозавад из Гедеры.
1CHR|12|6|Елузай, Иеримоф, Веалия, Шемария, Сафатия Харифиянин;
1CHR|12|7|Елкана, Ишшияху, Азариил, Иоезер и Иошавам, Кореяне;
1CHR|12|8|и Иоела и Зевадия, сыновья Иерохама, из Гедора.
1CHR|12|9|И из Гадитян перешли к Давиду в укрепление, в пустыню, люди мужественные, воинственные, вооруженные щитом и копьем; лица львиные – лица их, и они быстры как серны на горах.
1CHR|12|10|Главный Езер, второй Овадия, третий Елиав,
1CHR|12|11|четвертый Мишманна, пятый Иеремия,
1CHR|12|12|шестой Афай, седьмой Елиел,
1CHR|12|13|восьмой Иоханан, девятый Елзавад,
1CHR|12|14|десятый Иеремия, одиннадцатый Махбанай.
1CHR|12|15|Они из сыновей Гадовых [были] главами в войске: меньший над сотнею, и больший над тысячею.
1CHR|12|16|Они–то перешли Иордан в первый месяц, когда он выступает из берегов своих, и разогнали всех живших в долинах к востоку и западу.
1CHR|12|17|Пришли также и из сыновей Вениаминовых и Иудиных в укрепление к Давиду.
1CHR|12|18|Давид вышел навстречу им и сказал им: если с миром пришли вы ко мне, чтобы помогать мне, то да будет у меня с вами одно сердце; а если для того, чтобы коварно предать меня врагам моим, тогда как нет порока на руках моих, то да видит Бог отцов наших и рассудит.
1CHR|12|19|И объял дух Амасая, главу тридцати, [и сказал он]: мир тебе Давид, и с тобою, сын Иессеев; мир тебе, и мир помощникам твоим; ибо помогает тебе Бог твой. Тогда принял их Давид и поставил их во главе войска.
1CHR|12|20|И из колена Манассиина перешли [некоторые] к Давиду, когда он шел с Филистимлянами на войну против Саула, но не помогал им, потому что предводители Филистимские, посоветовавшись, отослали его, говоря: на нашу голову он перейдет к господину своему Саулу.
1CHR|12|21|Когда он возвращался в Секелаг, тогда перешли к нему из Манассиян: Аднах, Иозавад, Иедиаел, Михаил, Иозавад, Елигу и Цилльфай, тысяченачальники у Манассиян.
1CHR|12|22|И они помогали Давиду против полчищ, ибо все это были люди храбрые и были начальниками в войске.
1CHR|12|23|Так с каждым днем приходили к Давиду на помощь до того, что его ополчение стало велико, как ополчение Божие.
1CHR|12|24|Вот число главных в войске, которые пришли к Давиду в Хеврон, чтобы передать ему царство Саулово, по слову Господню:
1CHR|12|25|сыновей Иудиных, носящих щит и копье, было шесть тысяч восемьсот готовых к войне;
1CHR|12|26|из сыновей Симеоновых, людей храбрых, в войске было семь тысяч и сто;
1CHR|12|27|из сыновей Левииных четыре тысячи шестьсот;
1CHR|12|28|и Иоддай, князь от [племени] Аарона, и с ним три тысячи семьсот;
1CHR|12|29|и Садок, мужественный юноша, и род его, двадцать два начальника;
1CHR|12|30|из сыновей Вениаминовых, братьев Сауловых, три тысячи, – но еще многие из них держались дома Саулова;
1CHR|12|31|из сыновей Ефремовых двадцать тысяч восемьсот людей мужественных, людей именитых в родах своих;
1CHR|12|32|из полуколена Манассиина восемнадцать тысяч, которые вызваны были поименно, чтобы пойти воцарить Давида;
1CHR|12|33|из сынов Иссахаровых [пришли] люди разумные, которые знали, что когда надлежало делать Израилю, – их было двести главных, и все братья их следовали слову их;
1CHR|12|34|из [колена] Завулонова готовых к сражению, вооруженных всякими военными оружиями, пятьдесят тысяч, в строю, единодушных;
1CHR|12|35|из [колена] Неффалимова тысяча вождей и с ними тридцать семь тысяч с щитами и копьями;
1CHR|12|36|из [колена] Данова готовых к войне двадцать восемь тысяч шестьсот;
1CHR|12|37|от Асира воинов, готовых к сражению, сорок тысяч;
1CHR|12|38|из–за Иордана, от колена Рувимова, Гадова и полуколена Манассиина, сто двадцать тысяч, со всяким воинским оружием.
1CHR|12|39|Все эти воины, в строю, от полного сердца пришли в Хеврон воцарить Давида над всем Израилем. Да и все прочие Израильтяне были единодушны, чтобы воцарить Давида.
1CHR|12|40|И пробыли там у Давида три дня, ели и пили, потому что братья их [все] приготовили для них;
1CHR|12|41|да и близкие к ним, даже до [колена] Иссахарова, Завулонова и Неффалимова, привозили все съестное на ослах, и верблюдах, и мулах, и волах: муку, смоквы, и изюм, и вино, и елей, и крупного и мелкого скота множество, так как радость была для Израиля.
1CHR|13|1|И советовался Давид с тысяченачальниками, сотниками и со всеми вождями,
1CHR|13|2|и сказал [Давид] всему собранию Израильтян: если угодно вам, и если на то будет воля Господа Бога нашего, пошлем повсюду к прочим братьям нашим, по всей земле Израильской, и вместе с ними к священникам и левитам, в города и селения их, чтобы они собрались к нам;
1CHR|13|3|и перенесем к себе ковчег Бога нашего, потому что во дни Саула мы не обращались к нему.
1CHR|13|4|И сказало все собрание: "да будет так", потому что это дело всему народу казалось справедливым.
1CHR|13|5|Так собрал Давид всех Израильтян, от Шихора Египетского до входа в Емаф, чтобы перенести ковчег Божий из Кириаф–Иарима.
1CHR|13|6|И пошел Давид и весь Израиль в Кириаф–Иарим, что в Иудее, чтобы перенести оттуда ковчег Бога, Господа, седящего на Херувимах, на котором нарицается имя [Его].
1CHR|13|7|И повезли ковчег Божий на новой колеснице из дома Авинадава; и Оза и Ахия вели колесницу.
1CHR|13|8|Давид же и все Израильтяне играли пред Богом из всей силы, с пением, на цитрах и псалтирях, и тимпанах, и кимвалах и трубах.
1CHR|13|9|Когда дошли до гумна Хидона, Оза простер руку свою, чтобы придержать ковчег, ибо волы наклонили его.
1CHR|13|10|Но Господь разгневался на Озу, и поразил его за то, что он простер руку свою к ковчегу; и он умер тут же пред лицем Божиим.
1CHR|13|11|И опечалился Давид, что Господь поразил Озу. И назвал то место поражением Озы; так называется оно и до сего дня.
1CHR|13|12|И устрашился Давид Бога в день тот, и сказал: как я внесу к себе ковчег Божий?
1CHR|13|13|И не повез Давид ковчега к себе, в город Давидов, а обратил его к дому Аведдара Гефянина.
1CHR|13|14|И оставался ковчег Божий у Аведдара, в доме его, три месяца, и благословил Господь дом Аведдара и все, что у него.
1CHR|14|1|И послал Хирам, царь Тирский, к Давиду послов, и кедровые деревья, и каменщиков, и плотников, чтобы построить ему дом.
1CHR|14|2|Когда узнал Давид, что утвердил его Господь царем над Израилем, что вознесено высоко царство его, ради народа его Израиля,
1CHR|14|3|тогда взял Давид еще жен в Иерусалиме, и родил Давид еще сыновей и дочерей.
1CHR|14|4|И вот имена родившихся у него в Иерусалиме: Самус, Совав, Нафан, Соломон,
1CHR|14|5|Евеар, Елисуа, Елфалет,
1CHR|14|6|Ногах, Нафек, Иафиа,
1CHR|14|7|и Елисама, Веелиада и Елифалеф.
1CHR|14|8|И услышали Филистимляне, что помазан Давид в царя над всем Израилем, и поднялись все Филистимляне искать Давида. И услышал Давид [об] [этом] и пошел против них.
1CHR|14|9|И Филистимляне пришли и расположились в долине Рефаимов.
1CHR|14|10|И вопросил Давид Бога, говоря: идти ли мне против Филистимлян, и предашь ли их в руки мои? И сказал ему Господь: иди, и Я предам их в руки твои.
1CHR|14|11|И пошли они в Ваал–Перацим, и поразил их там Давид; и сказал Давид: сломил Бог врагов моих рукою моею, как прорыв воды. Посему и дали имя месту тому: Ваал–Перацим.
1CHR|14|12|И оставили там [Филистимляне] богов своих, и повелел Давид, и сожжены они огнем.
1CHR|14|13|И [пришли] опять Филистимляне и расположились по долине.
1CHR|14|14|И еще вопросил Давид Бога, и сказал ему Бог: не ходи [прямо] на них, уклонись от них и иди к ним со стороны тутовых дерев;
1CHR|14|15|и когда услышишь шум как бы шагов на вершинах тутовых дерев, тогда вступи в битву, ибо вышел Бог пред тобою, чтобы поразить стан Филистимлян.
1CHR|14|16|И сделал Давид, как повелел ему Бог; и поразили стан Филистимский, от Гаваона до Газера.
1CHR|14|17|И пронеслось имя Давидово по всем землям, и Господь сделал его страшным для всех народов.
1CHR|15|1|И построил он себе домы в городе Давидовом, и приготовил место для ковчега Божия, и устроил для него скинию.
1CHR|15|2|Тогда сказал Давид: [никто] не должен носить ковчега Божия, кроме левитов, потому что их избрал Господь на то, чтобы носить ковчег Божий и служить Ему во веки.
1CHR|15|3|И собрал Давид всех Израильтян в Иерусалим, чтобы внести ковчег Господень на место его, которое он для него приготовил.
1CHR|15|4|И созвал Давид сыновей Аароновых и левитов:
1CHR|15|5|из сыновей Каафовых, Уриила начальника и братьев его – сто двадцать [человек];
1CHR|15|6|из сыновей Мерариных, Асаию начальника и братьев его – двести двадцать [человек];
1CHR|15|7|из сыновей Гирсоновых, Иоиля начальника и братьев его – сто тридцать [человек];
1CHR|15|8|из сыновей Елисафановых, Шемаию начальника и братьев его – двести;
1CHR|15|9|из сыновей Хевроновых, Елиела начальника и братьев его – восемьдесят;
1CHR|15|10|из сыновей Уззииловых, Аминадава начальника и братьев его – сто двенадцать.
1CHR|15|11|И призвал Давид священников: Садока и Авиафара, и левитов: Уриила, Асаию, Иоиля, Шемаию, Елиела и Аминадава,
1CHR|15|12|и сказал им: вы, начальники родов левитских, освятитесь сами и братья ваши, и принесите ковчег Господа Бога Израилева на [место], [которое] я приготовил для него;
1CHR|15|13|ибо как прежде не вы это [делали], то Господь Бог наш поразил нас за то, что мы не взыскали Его, как должно.
1CHR|15|14|И освятились священники и левиты для того, чтобы нести ковчег Господа, Бога Израилева.
1CHR|15|15|И понесли сыновья левитов ковчег Божий, как заповедал Моисей по слову Господа, на плечах, на шестах.
1CHR|15|16|И приказал Давид начальникам левитов поставить братьев своих певцов с музыкальными орудиями, с псалтирями и цитрами и кимвалами, чтобы они громко возвещали глас радования.
1CHR|15|17|И поставили левиты Емана, сына Иоилева, и из братьев его, Асафа, сына Верехиина, а из сыновей Мерариных, братьев их, Ефана, сына Кушаии;
1CHR|15|18|и с ними братьев их второстепенных: Захарию, Бена, Иаазиила, Шемирамофа, Иехиила, Унния, Елиава, Ванею, Маасея, Маттафию, Елифлеуя, Микнея и Овед–Едома и Иеиела, привратников.
1CHR|15|19|Еман, Асаф и Ефан играли громко на медных кимвалах,
1CHR|15|20|а Захария, Азиил, Шемирамоф, Иехиил, Унний, Елиав, Маасей и Ванея – на псалтирях, тонким голосом.
1CHR|15|21|Маттафия же, Елифлеуй, Микней, Овед–Едом, Иеиел и Азазия – на цитрах, чтобы делать начало.
1CHR|15|22|А Хенания, начальник левитов, был учитель пения, потому что был искусен в нем.
1CHR|15|23|Верехия и Елкана были придверниками у ковчега.
1CHR|15|24|Шевания, Иосафат, Нафанаил, Амасай, Захария, Ванея и Елиезер, священники, трубили трубами пред ковчегом Божиим. Овед–Едом и Иехия [были] придверниками у ковчега.
1CHR|15|25|Так Давид и старейшины Израилевы и тысяченачальники пошли перенести ковчег завета Господня из дома Овед–Едомова с веселием.
1CHR|15|26|И когда Бог помог левитам, несшим ковчег завета Господня, тогда закололи в жертву семь тельцов и семь овнов.
1CHR|15|27|Давид был одет в виссонную одежду, [а также] и все левиты, несшие ковчег, и певцы, и Хенания начальник музыкантов и певцов. На Давиде же был [еще] льняной ефод.
1CHR|15|28|Так весь Израиль вносил ковчег завета Господня с восклицанием, при звуке рога и труб и кимвалов, играя на псалтирях и цитрах.
1CHR|15|29|Когда ковчег завета Господня входил в город Давидов, Мелхола, дочь Саулова, смотрела в окно и, увидев царя Давида, скачущего и веселящегося, уничижила его в сердце своем.
1CHR|16|1|И принесли ковчег Божий, и поставили его среди скинии, которую устроил для него Давид, и вознесли Богу всесожжения и мирные жертвы.
1CHR|16|2|Когда Давид окончил всесожжения и приношение мирных жертв, то благословил народ именем Господа
1CHR|16|3|и роздал всем Израильтянам, и мужчинам и женщинам, по одному хлебу и по куску мяса и по кружке вина,
1CHR|16|4|и поставил на службу пред ковчегом Господним [некоторых] из левитов, чтобы они славословили, благодарили и превозносили Господа Бога Израилева:
1CHR|16|5|Асафа главным, вторым по нем Захарию, Иеиела, Шемирамофа, Иехиила, Маттафию, Елиава, и Ванею, Овед–Едома и Иеиела с псалтирями и цитрами, и Асафа для игры на кимвалах,
1CHR|16|6|а Ванею и Озиила, священников, [чтобы] постоянно [трубили] пред ковчегом завета Божия.
1CHR|16|7|В этот день Давид в первый раз дал псалом для славословия Господу чрез Асафа и братьев его:
1CHR|16|8|славьте Господа, провозглашайте имя Его; возвещайте в народах дела Его;
1CHR|16|9|пойте Ему, бряцайте Ему; поведайте о всех чудесах Его;
1CHR|16|10|хвалитесь именем Его святым; да веселится сердце ищущих Господа;
1CHR|16|11|взыщите Господа и силы Его, ищите непрестанно лица Его;
1CHR|16|12|поминайте чудеса, которые Он сотворил, знамения Его и суды уст Его,
1CHR|16|13|[вы], семя Израилево, рабы Его, сыны Иакова, избранные Его!
1CHR|16|14|Он Господь Бог наш; суды Его по всей земле.
1CHR|16|15|Помните вечно завет Его, слово, которое Он заповедал в тысячу родов,
1CHR|16|16|то, что завещал Аврааму, и в чем клялся Исааку,
1CHR|16|17|и что поставил Иакову в закон и Израилю в завет вечный,
1CHR|16|18|говоря: "тебе дам Я землю Ханаанскую, в наследственный удел вам".
1CHR|16|19|Они были тогда малочисленны и ничтожны, и пришельцы в ней,
1CHR|16|20|и переходили от народа к народу и из одного царства к другому народу;
1CHR|16|21|но Он никому не позволил обижать их, и обличал за них царей:
1CHR|16|22|"Не прикасайтеся к помазанным Моим, и пророкам Моим не делайте зла".
1CHR|16|23|Пойте Господу, вся земля, благовествуйте изо дня в день спасение Его.
1CHR|16|24|Возвещайте язычникам славу Его, всем народам чудеса Его,
1CHR|16|25|ибо велик Господь и достохвален, страшен паче всех богов.
1CHR|16|26|Ибо все боги народов ничто, а Господь небеса сотворил.
1CHR|16|27|Слава и величие пред лицем Его, могущество и радость на месте Его.
1CHR|16|28|Воздайте Господу, племена народов, воздайте Господу славу и честь,
1CHR|16|29|воздайте Господу славу имени Его. Возьмите дар, идите пред лице Его, поклонитесь Господу в благолепии святыни Его.
1CHR|16|30|Трепещи пред Ним, вся земля, ибо Он основал вселенную, она не поколеблется.
1CHR|16|31|Да веселятся небеса, да торжествует земля, и да скажут в народах: Господь царствует!
1CHR|16|32|Да плещет море и что наполняет его, да радуется поле и все, что на нем.
1CHR|16|33|Да ликуют вместе все дерева дубравные пред лицем Господа, ибо Он идет судить землю.
1CHR|16|34|Славьте Господа, ибо вовек милость Его,
1CHR|16|35|и скажите: спаси нас, Боже, Спаситель наш! Собери нас и избавь нас от народов, да славим святое имя Твое и да хвалимся славою Твоею!
1CHR|16|36|Благословен Господь Бог Израилев, от века и до века! И сказал весь народ: аминь! аллилуия!
1CHR|16|37|Давид оставил там, пред ковчегом завета Господня, Асафа и братьев его, чтоб они служили пред ковчегом постоянно, каждый день,
1CHR|16|38|и Овед–Едома и братьев его, шестьдесят восемь [человек]; Овед–Едома, сына Идифунова, и Хосу – привратниками,
1CHR|16|39|а Садока священника и братьев его священников пред жилищем Господним, что на высоте в Гаваоне,
1CHR|16|40|для возношения всесожжений Господу на жертвеннике всесожжения постоянно, утром и вечером, и для всего, что написано в законе Господа, который Он заповедал Израилю;
1CHR|16|41|и с ними Емана и Идифуна и прочих избранных, которые назначены поименно, чтобы славить Господа, ибо навек милость Его.
1CHR|16|42|При них Еман и Идифун прославляли Бога, играя на трубах, кимвалах и разных музыкальных орудиях; сыновей же Идифуна [поставил] при вратах.
1CHR|16|43|И пошел весь народ, каждый в свой дом; возвратился и Давид, чтобы благословить дом свой.
1CHR|17|1|Когда Давид жил в доме своем, то сказал Давид Нафану пророку: вот, я живу в доме кедровом, а ковчег завета Господня под шатром.
1CHR|17|2|И сказал Нафан Давиду: все, что у тебя на сердце, делай, ибо с тобою Бог.
1CHR|17|3|Но в ту же ночь было слово Божие к Нафану:
1CHR|17|4|пойди и скажи рабу Моему Давиду: так говорит Господь: не ты построишь Мне дом для обитания,
1CHR|17|5|ибо Я не жил в доме с того дня, как вывел сынов Израиля, и до сего дня, а [ходил] из скинии в скинию и из жилища [в жилище].
1CHR|17|6|Где ни ходил Я со всем Израилем, сказал ли Я хотя слово которому–либо из судей Израильских, которым Я повелел пасти народ Мой: зачем вы не построите Мне дома кедрового?
1CHR|17|7|И теперь так скажи рабу Моему Давиду: так говорит Господь Саваоф: Я взял тебя от стада овец, чтобы ты был вождем народа Моего Израиля;
1CHR|17|8|и был с тобою везде, куда ты ни ходил, и истребил всех врагов твоих пред лицем твоим, и сделал имя твое, как имя великих на земле;
1CHR|17|9|и Я устроил место для народа Моего Израиля, и укоренил его, и будет он спокойно жить на месте своем, и не будет более тревожим, и нечестивые не станут больше теснить его, как прежде,
1CHR|17|10|в те дни, когда Я поставил судей над народом Моим Израилем, и Я смирил всех врагов твоих, и возвещаю тебе, что Господь устроит тебе дом.
1CHR|17|11|Когда исполнятся дни твои, и ты отойдешь к отцам твоим, тогда Я восставлю семя твое после тебя, которое будет из сынов твоих, и утвержу царство его.
1CHR|17|12|Он построит Мне дом, и утвержу престол его на веки.
1CHR|17|13|Я буду ему отцом, и он будет Мне сыном, – и милости Моей не отниму от него, как Я отнял от того, который был прежде тебя.
1CHR|17|14|Я поставлю его в доме Моем и в царстве Моем на веки, и престол его будет тверд вечно.
1CHR|17|15|Все эти слова и все видение точно пересказал Нафан Давиду.
1CHR|17|16|И пришел царь Давид, и стал пред лицем Господним, и сказал: кто я, Господи Боже, и что такое дом мой, что Ты так возвысил меня?
1CHR|17|17|Но и этого еще мало показалось в очах Твоих, Боже; Ты возвещаешь о доме раба Твоего вдаль, и взираешь на меня, как на человека великого, Господи Боже!
1CHR|17|18|Что еще может прибавить пред Тобою Давид для возвеличения раба Твоего? Ты знаешь раба Твоего!
1CHR|17|19|Господи! для раба Твоего, по сердцу Твоему, Ты делаешь все это великое, чтобы явить всякое величие.
1CHR|17|20|Господи! Нет подобного Тебе, и нет Бога, кроме Тебя, по всему, что слышали мы своими ушами.
1CHR|17|21|И кто подобен народу Твоему Израилю, единственному народу на земле, к которому приходил Бог, [чтоб] искупить его Себе в народ, сделать Себе имя великим и страшным делом – прогнанием народов от лица народа Твоего, который Ты избавил из Египта.
1CHR|17|22|Ты соделал народ Твой Израиля Своим собственным народом навек, и Ты, Господи, стал Богом его.
1CHR|17|23|Итак теперь, о, Господи, слово, которое Ты сказал о рабе Твоем и о доме его, утверди навек, и сделай, как Ты сказал.
1CHR|17|24|И да пребудет и возвеличится имя Твое во веки, чтобы говорили: Господь Саваоф, Бог Израилев, есть Бог над Израилем, и дом раба Твоего Давида да будет тверд пред лицем Твоим.
1CHR|17|25|Ибо Ты, Боже мой, открыл рабу Твоему, что Ты устроишь ему дом, поэтому раб Твой и дерзнул молиться пред Тобою.
1CHR|17|26|И ныне, Господи, Ты Бог, и Ты сказал о рабе Твоем такое благо.
1CHR|17|27|Начни же благословлять дом раба Твоего, чтоб он был вечно пред лицем Твоим. Ибо если Ты, Господи, благословишь, то будет он благословен вовек.
1CHR|18|1|После сего Давид поразил Филистимлян и смирил их, и взял Геф и зависящие от него города из руки Филистимлян.
1CHR|18|2|Он поразил также Моавитян, – и сделались Моавитяне рабами Давида, принося ему дань.
1CHR|18|3|И поразил Давид Адраазара, царя Сувского, в Емафе, когда тот шел утвердить власть свою при реке Евфрате.
1CHR|18|4|И взял Давид у него тысячу колесниц, семь тысяч всадников и двадцать тысяч пеших, и разрушил Давид все колесницы, оставив из них [только] сто.
1CHR|18|5|Сирияне Дамасские пришли было на помощь к Адраазару, царю Сувскому, но Давид поразил двадцать две тысячи Сириян.
1CHR|18|6|И поставил Давид [охранное войско] в Сирии Дамасской, и сделались Сирияне рабами Давида, принося ему дань. И помогал Господь Давиду везде, куда он ни ходил.
1CHR|18|7|И взял Давид золотые щиты, которые были у рабов Адраазара, и принес их в Иерусалим.
1CHR|18|8|А из Тивхавы и Куна, городов Адраазаровых, взял Давид весьма много меди. Из нее Соломон сделал медное море и столбы и медные сосуды.
1CHR|18|9|И услышал Фой, царь Имафа, что Давид поразил все войско Адраазара, царя Сувского.
1CHR|18|10|И послал Иорама, сына своего, к царю Давиду, приветствовать его и благодарить за то, что он воевал с Адраазаром и поразил его, ибо Фой был в войне с Адраазаром, – и [с ним] всякие сосуды золотые, серебряные и медные.
1CHR|18|11|И посвятил их царь Давид Господу вместе с серебром и золотом, которое он взял от всех народов: от Идумеян, Моавитян, Аммонитян, Филистимлян и от Амаликитян.
1CHR|18|12|И Авесса, сын Саруи, поразил Идумеян на долине Соляной восемнадцать тысяч;
1CHR|18|13|и поставил в Идумее охранное войско, и сделались все Идумеяне рабами Давиду. Господь помогал Давиду везде, куда он ни ходил.
1CHR|18|14|И царствовал Давид над всем Израилем, и творил суд и правду всему народу своему.
1CHR|18|15|Иоав, сын Саруи, [был] начальником войска, Иосафат, сын Ахилуда, дееписателем,
1CHR|18|16|Садок, сын Ахитува, и Авимелех, сын Авиафара, священниками, а Суса писцом,
1CHR|18|17|Ванея, сын Иодая, над Хелефеями и Фелефеями, а сыновья Давидовы – первыми при царе.
1CHR|19|1|После сего умер Наас, царь Аммонитский, и воцарился сын его вместо него.
1CHR|19|2|И сказал Давид: окажу я милость Аннону, сыну Наасову, за благодеяние, которое отец его оказал мне. И послал Давид послов утешить его об отце его; и пришли слуги Давидовы в землю Аммонитскую, к Аннону, чтобы утешить его.
1CHR|19|3|Но князья Аммонитские сказали Аннону: неужели ты думаешь, что Давид из уважения к отцу твоему прислал к тебе утешителей? Не для того ли пришли слуги его к тебе, чтобы разведать и высмотреть землю и разорить ее?
1CHR|19|4|И взял Аннон слуг Давидовых и обрил их, и обрезал одежды их наполовину до чресл и отпустил их.
1CHR|19|5|И пошли они. И донесено было Давиду о людях сих, и он послал им навстречу, так как они были очень обесчещены; и сказал царь: останьтесь в Иерихоне, пока отрастут бороды ваши, и тогда возвратитесь.
1CHR|19|6|Когда Аммонитяне увидели, что они сделались ненавистными Давиду, тогда послал Аннон и Аммонитяне тысячу талантов серебра, чтобы нанять себе колесниц и всадников из Сирии Месопотамской и из Сирии Мааха и из Сувы.
1CHR|19|7|И наняли себе тридцать две тысячи колесниц и царя Мааха с народом его, которые пришли и расположились станом пред Медевою. И Аммонитяне собрались из городов своих и выступили на войну.
1CHR|19|8|Когда услышал об этом Давид, то послал Иоава со всем войском храбрых.
1CHR|19|9|И выступили Аммонитяне и выстроились к сражению у ворот города, а цари, которые пришли, отдельно в поле.
1CHR|19|10|Иоав, видя, что предстоит ему сражение спереди и сзади, избрал воинов из всех отборных в Израиле и выстроил [их] против Сириян.
1CHR|19|11|А остальную часть народа поручил Авессе, брату своему, чтоб они выстроились против Аммонитян.
1CHR|19|12|И сказал он: если Сирияне будут одолевать меня, то ты поможешь мне, а если Аммонитяне будут одолевать тебя, то я помогу тебе.
1CHR|19|13|Будь мужествен, и будем твердо стоять за народ наш и за города Бога нашего, – и Господь пусть сделает, что ему угодно.
1CHR|19|14|И вступил Иоав и люди, которые были у него, в сражение с Сириянами, и они побежали от него.
1CHR|19|15|Аммонитяне же, увидев, что Сирияне бегут, и сами побежали от Авессы, брата его, и ушли в город. И пришел Иоав в Иерусалим.
1CHR|19|16|Сирияне, видя, что они поражены Израильтянами, отправили послов и вывели Сириян, которые были по ту сторону реки, и Совак, военачальник Адраазаров, предводительствовал ими.
1CHR|19|17|Когда донесли об этом Давиду, он собрал всех Израильтян, перешел Иордан и, придя к ним, выстроился против них; и вступил Давид в сражение с Сириянами, и они сразились с ним.
1CHR|19|18|И Сирияне побежали от Израильтян, и истребил Давид у Сириян семь тысяч колесниц и сорок тысяч пеших, и Совака военачальника умертвил.
1CHR|19|19|Когда увидели слуги Адраазара, что они поражены Израильтянами, заключили с Давидом мир и подчинились ему. И не хотели Сирияне помогать более Аммонитянам.
1CHR|20|1|Через год, в то время когда цари выходят [на войну], вывел Иоав войско и стал разорять землю Аммонитян, и пришел и осадил Равву. Давид же оставался в Иерусалиме. Иоав, завоевав Равву, разрушил ее.
1CHR|20|2|И взял Давид венец царя их с головы его, и в нем оказалось весу талант золота, и драгоценные камни были на нем; и был он возложен на голову Давида. И добычи очень много вынес из города.
1CHR|20|3|А народ, который был в нем, вывел и умерщвлял их пилами, железными молотилами и секирами. Так поступил Давид со всеми городами Аммонитян, и возвратился Давид и весь народ в Иерусалим.
1CHR|20|4|После того началась война с Филистимлянами в Газере. Тогда Совохай Хушатянин поразил Сафа, одного из потомков Рефаимов. И они усмирились.
1CHR|20|5|И опять была война с Филистимлянами. Тогда Елханам, сын Иаира, поразил Лахмия, брата Голиафова, Гефянина, у которого древко копья было, как навой у ткачей.
1CHR|20|6|Было еще сражение в Гефе. Там был один рослый человек, у которого было по шести пальцев, [всего] двадцать четыре. И он также был из потомков Рефаимов.
1CHR|20|7|Он поносил Израиля, но Ионафан, сын Шимы, брата Давидова, поразил его.
1CHR|20|8|Это были родившиеся от Рефаимов в Гефе, и пали от руки Давида и от руки слуг его.
1CHR|21|1|И восстал сатана на Израиля, и возбудил Давида сделать счисление Израильтян.
1CHR|21|2|И сказал Давид Иоаву и начальствующим в народе: пойдите исчислите Израильтян, от Вирсавии до Дана, и представьте мне, чтоб я знал число их.
1CHR|21|3|И сказал Иоав: да умножит Господь народ Свой во сто раз против того, сколько есть его. Не все ли они, господин мой царь, рабы господина моего? Для чего же требует сего господин мой? Чтобы вменилось это в вину Израилю?
1CHR|21|4|Но царское слово превозмогло Иоава; и пошел Иоав, и обошел всего Израиля, и пришел в Иерусалим.
1CHR|21|5|И подал Иоав Давиду список народной переписи, и было всех Израильтян тысяча тысяч, и сто тысяч мужей, обнажающих меч, и Иудеев – четыреста семьдесят тысяч, обнажающих меч.
1CHR|21|6|А левитов и Вениаминян он не исчислял между ними, потому что царское слово противно было Иоаву.
1CHR|21|7|И не угодно было в очах Божиих дело сие, и Он поразил Израиля.
1CHR|21|8|И сказал Давид Богу: весьма согрешил я, что сделал это. И ныне прости вину раба Твоего, ибо я поступил очень безрассудно.
1CHR|21|9|И говорил Господь Гаду, прозорливцу Давидову, и сказал:
1CHR|21|10|пойди и скажи Давиду: так говорит Господь: три [наказания] Я предлагаю тебе, избери себе одно из них, – и Я пошлю его на тебя.
1CHR|21|11|И пришел Гад к Давиду и сказал ему: так говорит Господь: избирай себе:
1CHR|21|12|или три года – голод, или три месяца будешь ты преследуем неприятелями твоими и меч врагов твоих будет досягать [до тебя]; или три дня – меч Господень и язва на земле и Ангел Господень, истребляющий во всех пределах Израиля. Итак, рассмотри, что мне отвечать Пославшему меня с словом.
1CHR|21|13|И сказал Давид Гаду: тяжело мне очень, но пусть лучше впаду в руки Господа, ибо весьма велико милосердие Его, только бы не впасть мне в руки человеческие.
1CHR|21|14|И послал Господь язву на Израиля, и умерло Израильтян семьдесят тысяч человек.
1CHR|21|15|И послал Бог Ангела в Иерусалим, чтобы истреблять его. И когда он начал истреблять, увидел Господь и пожалел о сем бедствии, и сказал Ангелу–истребителю: довольно! теперь опусти руку твою. Ангел же Господень стоял [тогда] над гумном Орны Иевусеянина.
1CHR|21|16|И поднял Давид глаза свои, и увидел Ангела Господня, стоящего между землею и небом, с обнаженным в руке его мечом, простертым на Иерусалим; и пал Давид и старейшины, покрытые вретищем, на лица свои.
1CHR|21|17|И сказал Давид Богу: не я ли велел исчислить народ? я согрешил, я сделал зло, а эти овцы что сделали? Господи, Боже мой! да будет рука Твоя на мне и на доме отца моего, а не на народе Твоем, чтобы погубить [его].
1CHR|21|18|И Ангел Господень сказал Гаду, чтобы тот сказал Давиду: пусть Давид придет и поставит жертвенник Господу на гумне Орны Иевусеянина.
1CHR|21|19|И пошел Давид, по слову Гада, которое он говорил именем Господним.
1CHR|21|20|Орна обратился, увидел Ангела, и четыре сына его с ним скрылись. Орна молотил тогда пшеницу.
1CHR|21|21|И пришел Давид к Орне. Орна, взглянув и увидев Давида, вышел из гумна и поклонился Давиду лицем до земли.
1CHR|21|22|И сказал Давид Орне: отдай мне место под гумном, я построю на нем жертвенник Господу; за настоящую цену отдай мне его, чтобы прекратилось истребление народа.
1CHR|21|23|И сказал Орна Давиду: возьми себе; пусть делает господин мой царь что ему угодно; вот я отдаю и волов на всесожжение, и молотильные орудия на дрова, и пшеницу на приношение; все это отдаю даром.
1CHR|21|24|И сказал царь Давид Орне: нет, я хочу купить у тебя за настоящую цену, ибо не стану я приносить твоей собственности Господу, и не буду приносить во всесожжение [взятого] даром.
1CHR|21|25|И дал Давид Орне за это место шестьсот сиклей золота.
1CHR|21|26|И соорудил там Давид жертвенник Господу и вознес всесожжения и мирные жертвы; и призвал Господа, и Он услышал его, [послав] огонь с неба на жертвенник всесожжения.
1CHR|21|27|И сказал Господь Ангелу: возврати меч твой в ножны его.
1CHR|21|28|В это время Давид, видя, что Господь услышал его на гумне Орны Иевусеянина, принес там жертву.
1CHR|21|29|Скиния же Господня, которую сделал Моисей в пустыне, и жертвенник всесожжения [находились] в то время на высоте в Гаваоне.
1CHR|21|30|И не мог Давид пойти туда, чтобы взыскать Бога, потому что устрашен был мечом Ангела Господня.
1CHR|22|1|И сказал Давид: вот дом Господа Бога и вот жертвенник для всесожжений Израиля.
1CHR|22|2|И приказал Давид собрать пришельцев, находившихся в земле Израильской, и поставил каменотесов, чтобы обтесывать камни для построения дома Божия.
1CHR|22|3|И множество железа для гвоздей к дверям ворот и для связей заготовил Давид, и множество меди без весу,
1CHR|22|4|и кедровых дерев без счету, потому что Сидоняне и Тиряне доставили Давиду множество кедровых дерев.
1CHR|22|5|И сказал Давид: Соломон, сын мой, молод и малосилен, а дом, который следует выстроить для Господа, должен быть весьма величествен, на славу и украшение пред всеми землями: итак буду я заготовлять для него. И заготовил Давид до смерти своей много.
1CHR|22|6|И призвал Соломона, сына своего, и завещал ему построить дом Господу Богу Израилеву.
1CHR|22|7|И сказал Давид Соломону: сын мой! у меня было на сердце построить дом во имя Господа, Бога моего,
1CHR|22|8|но было ко мне слово Господне, и сказано: "ты пролил много крови и вел большие войны; ты не должен строить дома имени Моему, потому что пролил много крови на землю пред лицем Моим.
1CHR|22|9|Вот, у тебя родится сын: он будет человек мирный; Я дам ему покой от всех врагов его кругом: посему имя ему будет Соломон. И мир и покой дам Израилю во дни его.
1CHR|22|10|Он построит дом имени Моему, и он будет Мне сыном, а Я ему отцом, и утвержу престол царства его над Израилем навек".
1CHR|22|11|И ныне, сын мой! да будет Господь с тобою, чтобы ты был благоуспешен и построил дом Господу Богу твоему, как Он говорил о тебе.
1CHR|22|12|Да даст тебе Господь смысл и разум, и поставит тебя над Израилем; и соблюди закон Господа Бога твоего.
1CHR|22|13|Тогда ты будешь благоуспешен, если будешь стараться исполнять уставы и законы, которые заповедал Господь Моисею для Израиля. Будь тверд и мужествен, не бойся и не унывай.
1CHR|22|14|И вот, я при скудости моей приготовил для дома Господня сто тысяч талантов золота и тысячу тысяч талантов серебра, а меди и железу нет веса, потому что их множество; и дерева и камни я также заготовил, а ты еще прибавь к этому.
1CHR|22|15|У тебя множество рабочих, и каменотесов, резчиков и плотников, и всяких способных на всякое дело;
1CHR|22|16|золоту, серебру и меди и железу нет счета: начни и делай; Господь будет с тобою.
1CHR|22|17|И завещал Давид всем князьям Израилевым помогать Соломону, сыну его:
1CHR|22|18|не с вами ли Господь Бог наш, давший вам покой со всех сторон? потому что Он предал в руки мои жителей земли, и покорилась земля пред Господом и пред народом Его.
1CHR|22|19|Итак расположите сердце ваше и душу вашу к тому, чтобы взыскать Господа Бога вашего. Встаньте и постройте святилище Господу Богу, чтобы перенести ковчег завета Господня и священные сосуды Божии в дом, созидаемый имени Господню.
1CHR|23|1|Давид, состарившись и насытившись [жизнью], воцарил над Израилем сына своего Соломона.
1CHR|23|2|И собрал всех князей Израилевых и священников и левитов,
1CHR|23|3|и исчислены были левиты, от тридцати лет и выше, и было число их, считая поголовно, тридцать восемь тысяч человек.
1CHR|23|4|Из них [назначены] для дела в доме Господнем двадцать четыре тысячи, писцов же и судей шесть тысяч,
1CHR|23|5|и четыре тысячи привратников, и четыре тысячи прославляющих Господа на [музыкальных] орудиях, которые он сделал для прославления.
1CHR|23|6|И разделил их Давид на череды по сынам Левия – Гирсону, Каафу и Мерари.
1CHR|23|7|Из Гирсонян – Лаедан и Шимей.
1CHR|23|8|Сыновья Лаедана: первый Иехиил, Зефам и Иоиль, трое.
1CHR|23|9|Сыновья Шимея: Шеломиф, Хазиил и Гаран, трое. Они главы поколений Лаедановых.
1CHR|23|10|Еще сыновья Шимея: Иахаф, Зиза, Иеуш и Берия. Это сыновья Шимея, четверо.
1CHR|23|11|Иахаф был главным, Зиза вторым; Иеуш и Берия имели детей немного, и потому они были в одном счете при доме отца.
1CHR|23|12|Сыновья Каафа: Амрам, Ицгар, Хеврон и Озиил, четверо.
1CHR|23|13|Сыновья Амрама: Аарон и Моисей. Аарон отделен был на посвящение ко Святому Святых, он и сыновья его, на веки, чтобы совершать курение пред лицем Господа, чтобы служить Ему и благословлять именем Его на веки.
1CHR|23|14|А Моисей, человек Божий, [и] сыновья его причтены к колену Левиину.
1CHR|23|15|Сыновья Моисея: Гирсон и Елиезер.
1CHR|23|16|Сыновья Гирсона: первый был Шевуил.
1CHR|23|17|Сыновья Елиезера были: первый Рехавия. И не было у Елиезера других сыновей; у Рехавии же было очень много сыновей.
1CHR|23|18|Сыновья Ицгара: первый Шеломиф.
1CHR|23|19|Сыновья Хеврона: первый Иерия и второй Амария, третий Иахазиил и четвертый Иекамам.
1CHR|23|20|Сыновья Озиила: первый Миха и второй Ишшия.
1CHR|23|21|Сыновья Мерарины: Махли и Муши. Сыновья Махлия: Елеазар и Кис.
1CHR|23|22|И умер Елеазар, и не было у него сыновей, а только дочери; и взяли их за себя сыновья Киса, братья их.
1CHR|23|23|Сыновья Мушия: Махли, Едер и Иремоф – трое.
1CHR|23|24|Вот сыновья Левиины, по домам отцов их, главы семейств, по именному счислению их поголовно, которые отправляли дела служения в доме Господнем, от двадцати лет и выше.
1CHR|23|25|Ибо Давид сказал: Господь, Бог Израилев, дал покой народу Своему и водворил его в Иерусалиме на веки,
1CHR|23|26|и левитам не нужно носить скинию и всякие вещи ее для служения в ней.
1CHR|23|27|Посему, по последним повелениям Давида, исчислены левиты от двадцати лет и выше,
1CHR|23|28|чтоб они были при сынах Аароновых, для служения дому Господню, во дворе и в пристройках, для соблюдения чистоты всего святилища и для исполнения всякой службы при доме Божием,
1CHR|23|29|для наблюдения за хлебами предложения и пшеничною мукою для хлебного приношения и пресными лепешками, за печеным, жареным и за всякою мерою и весом,
1CHR|23|30|и чтобы становились каждое утро благодарить и славословить Господа, также и вечером,
1CHR|23|31|и при всех всесожжениях, возносимых Господу в субботы, в новомесячия и в праздники по числу, как предписано о них, – постоянно пред лицем Господа,
1CHR|23|32|и чтобы охраняли скинию откровения и святилище и сынов Аароновых, братьев своих, при службах дому Господню.
1CHR|24|1|И вот распределения сыновей Аароновых: сыновья Аарона: Надав, Авиуд, Елеазар и Ифамар.
1CHR|24|2|Надав и Авиуд умерли прежде отца своего, сыновей же не было у них, и потому священствовали Елеазар и Ифамар.
1CHR|24|3|И распределил их Давид – Садока из сыновей Елеазара, и Ахимелеха из сыновей Ифамара, поочередно на службу их.
1CHR|24|4|И нашлось, что между сынами Елеазара глав поколений более, нежели между сынами Ифамара. И он распределил их [так]: из сынов Елеазара шестнадцать глав семейств, а из сынов Ифамара восемь.
1CHR|24|5|Распределял же их по жребиям, потому что главными во святилище и главными пред Богом были из сынов Елеазара и из сынов Ифамара,
1CHR|24|6|и записывал их Шемаия, сын Нафанаила, писец из левитов, пред лицем царя и князей и пред священником Садоком и Ахимелехом, сыном Авиафара, и пред главами семейств священнических и левитских: брали [при] [бросании жребия] одно семейство из [рода] Елеазарова, потом брали из [рода] Ифамарова.
1CHR|24|7|И вышел первый жребий Иегоиариву, второй Иедаии,
1CHR|24|8|третий Хариму, четвертый Сеориму,
1CHR|24|9|пятый Малхию, шестой Миямину,
1CHR|24|10|седьмой Гаккоцу, восьмой Авии,
1CHR|24|11|девятый Иешую, десятый Шехании,
1CHR|24|12|одиннадцатый Елиашиву, двенадцатый Иакиму,
1CHR|24|13|тринадцатый Хушаю, четырнадцатый Иешеваву,
1CHR|24|14|пятнадцатый Вилге, шестнадцатый Имеру,
1CHR|24|15|семнадцатый Хезиру, восемнадцатый Гапицецу,
1CHR|24|16|девятнадцатый Петахии, двадцатый Иезекиилю,
1CHR|24|17|двадцать первый Иахину, двадцать второй Гамулу,
1CHR|24|18|двадцать третий Делаии, двадцать четвертый Маазии.
1CHR|24|19|Вот порядок их при служении их, как [им] приходить в дом Господень, по уставу их чрез Аарона, отца их, как заповедал ему Господь Бог Израилев.
1CHR|24|20|У прочих сыновей Левия – [распределение]: из сынов Амрама: Шуваил; из сынов Шуваила: Иедия;
1CHR|24|21|от Рехавии: из сынов Рехавии Ишшия был первый;
1CHR|24|22|от Ицгара: Шеломоф; из сыновей Шеломофа: Иахав;
1CHR|24|23|из сыновей [Хеврона]: первый Иерия, второй Амария, третий Иахазиил, четвертый Иекамам.
1CHR|24|24|[Из] сыновей Озиила: Миха; из сыновей Михи: Шамир.
1CHR|24|25|Брат Михи Ишшия; из сыновей Ишшии: Захария.
1CHR|24|26|Сыновья Мерари: Махли и Муши; [из] сыновей Иаазии: Бено.
1CHR|24|27|[Из] сыновей Мерари у Иаазии: Бено и Шогам, и Заккур и Иври.
1CHR|24|28|У Махлия – Елеазар; у него сыновей не было.
1CHR|24|29|У Киса: [из] сыновей Киса: Иерахмиил;
1CHR|24|30|сыновья Мушия: Махли, Едер и Иеримоф. Вот сыновья левитов по поколениям их.
1CHR|24|31|Бросали и они жребий, наравне с братьями своими, сыновьями Аароновыми, пред лицем царя Давида и Садока и Ахимелеха, и глав семейств священнических и левитских: глава семейства наравне с меньшим братом своим.
1CHR|25|1|И отделил Давид и начальники войска на службу сыновей Асафа, Емана и Идифуна, чтобы они провещавали на цитрах, псалтирях и кимвалах; и были отчислены они на дело служения своего:
1CHR|25|2|из сыновей Асафа: Заккур, Иосиф, Нефания и Ашарела сыновья Асафа, под руководством Асафа, игравшего по наставлению царя.
1CHR|25|3|От Идифуна сыновья Идифуна: Гедалия, Цери, Исаия, Семей, Хашавия и Маттафия, шестеро, под руководством отца своего Идифуна, игравшего на цитре во славу и хвалу Господа.
1CHR|25|4|От Емана сыновья Емана: Буккия, Матфания, Озиил, Шевуил и Иеримоф, Ханания, Ханани, Елиафа, Гиддалти, Ромамти–Езер, Иошбекаша, Маллофи, Гофир и Махазиоф.
1CHR|25|5|Все эти сыновья Емана, прозорливца царского, по словам Божиим, чтобы возвышать славу его. И дал Бог Еману четырнадцать сыновей и трех дочерей.
1CHR|25|6|Все они под руководством отца своего пели в доме Господнем с кимвалами, псалтирями и цитрами в служении в доме Божием, по указанию царя, или Асафа, Идифуна и Емана.
1CHR|25|7|И было число их с братьями их, обученными петь пред Господом, всех знающих [сие дело], двести восемьдесят восемь.
1CHR|25|8|И бросили они жребий о череде служения, малый наравне с большим, учители [наравне] с учениками.
1CHR|25|9|И вышел первый жребий Асафу, для Иосифа; второй Гедалии с братьями его и сыновьями его; их было двенадцать;
1CHR|25|10|третий Заккуру с сыновьями его и братьями его; их – двенадцать;
1CHR|25|11|четвертый Ицрию с сыновьями его и братьями его; их – двенадцать;
1CHR|25|12|пятый Нефании с сыновьями его и братьями его; их – двенадцать;
1CHR|25|13|шестой Буккии с сыновьями его и братьями его; их – двенадцать;
1CHR|25|14|седьмой Иесареле с сыновьями его и братьями его; их – двенадцать;
1CHR|25|15|восьмой Исаии с сыновьями его и братьями его; их – двенадцать;
1CHR|25|16|девятый Матфании с сыновьями его и братьями его; их – двенадцать;
1CHR|25|17|десятый Шимею с сыновьями его и братьями его; их – двенадцать;
1CHR|25|18|одиннадцатый Азариилу с сыновьями его и братьями его; их – двенадцать;
1CHR|25|19|двенадцатый Хашавии с сыновьями его и братьями его; их – двенадцать;
1CHR|25|20|тринадцатый Шуваилу с сыновьями его и братьями его; их – двенадцать;
1CHR|25|21|четырнадцатый Маттафии с сыновьями его и братьями его; их – двенадцать;
1CHR|25|22|пятнадцатый Иеримофу с сыновьями его и братьями его; их – двенадцать;
1CHR|25|23|шестнадцатый Ханании с сыновьями его и братьями его; их – двенадцать;
1CHR|25|24|семнадцатый Иошбекаше с сыновьями его и братьями его; их – двенадцать;
1CHR|25|25|восемнадцатый Ханани с сыновьями его и братьями его; их – двенадцать;
1CHR|25|26|девятнадцатый Маллофию с сыновьями его и братьями его; их – двенадцать;
1CHR|25|27|двадцатый Елиафе с сыновьями его и братьями его; их – двенадцать;
1CHR|25|28|двадцать первый Гофиру с сыновьями его и братьями его; их – двенадцать;
1CHR|25|29|двадцать второй Гиддалтию с сыновьями его и братьями его; их – двенадцать;
1CHR|25|30|двадцать третий Махазиофу с сыновьями его и братьями его; их – двенадцать;
1CHR|25|31|двадцать четвертый Ромамти–Езеру с сыновьями его и братьями его; их – двенадцать.
1CHR|26|1|Вот распределение привратников: из Кореян: Мешелемия, сын Корея, из сыновей Асафовых.
1CHR|26|2|Сыновья Мешелемии: первенец Захария, второй Иедиаил, третий Зевадия, четвертый Иафниил,
1CHR|26|3|пятый Елам, шестой Иегоханан, седьмой Елиегоэнай.
1CHR|26|4|Сыновья Овед–Едома: первенец Шемаия, второй Иегозавад, третий Иоах, четвертый Сахар, пятый Нафанаил,
1CHR|26|5|шестой Аммиил, седьмой Иссахар, восьмой Пеульфай, потому что Бог благословил его.
1CHR|26|6|У сына его Шемаии родились также сыновья, начальствовавшие в своем роде, потому что они были люди сильные.
1CHR|26|7|Сыновья Шемаии: Офни, Рефаил, Овед и Елзавад, братья его, люди сильные, Елия, Семахия.
1CHR|26|8|Все они из сыновей Овед–Едома; они и сыновья их, и братья их были люди прилежные и к службе способные: их было у Овед–Едома шестьдесят два.
1CHR|26|9|У Мешелемии сыновей и братьев, людей способных, [было] восемнадцать.
1CHR|26|10|У Хосы, из сыновей Мерариных, сыновья: Шимри главный, – хотя он не был первенцем, но отец его поставил его главным;
1CHR|26|11|второй Хелкия, третий Тевалия, четвертый Захария; всех сыновей и братьев у Хосы было тринадцать.
1CHR|26|12|Вот распределение привратников по главам семейств, способных на службу вместе с братьями их, для служения в доме Господнем.
1CHR|26|13|И бросили они жребии, как малый, так и большой, по своим семействам, на каждые ворота.
1CHR|26|14|И выпал жребий на восток Шелемии; и Захарии, сыну его, умному советнику, бросили жребий, и вышел ему жребий на север;
1CHR|26|15|Овед–Едому на юг, а сыновьям его при кладовых.
1CHR|26|16|Шупиму и Хосе на запад, у ворот Шаллехет, где дорога поднимается и где стража против стражи.
1CHR|26|17|К востоку по шести левитов, к северу по четыре, к югу по четыре, а у кладовых по два.
1CHR|26|18|К западу у притвора на дороге по четыре, а у самого притвора по два.
1CHR|26|19|Вот распределение привратников из сыновей Кореевых и сыновей Мерариных.
1CHR|26|20|Левиты же, братья их, [смотрели] за сокровищами дома Божия и за сокровищницами посвященных вещей.
1CHR|26|21|Сыновья Лаедана, сына Герсонова – от Лаедана, главы семейств от Лаедана Герсонского: Иехиел.
1CHR|26|22|Сыновья Иехиела: Зефам и Иоиль, брат его, [смотрели] за сокровищами дома Господня,
1CHR|26|23|вместе с потомками Амрама, Ицгара, Хеврона, Озиила.
1CHR|26|24|Шевуил, сын Гирсона, сына Моисеева, [был] главным смотрителем за сокровищницами.
1CHR|26|25|У брата его Елиезера сын Рехавия, у него сын Исаия, у него сын Иорам, у него сын Зихрий, у него сын Шеломиф.
1CHR|26|26|Шеломиф и братья его [смотрели] за всеми сокровищницами посвященных вещей, которые посвятил царь Давид и главы семейств и тысяченачальники, стоначальники и предводители войска.
1CHR|26|27|Из завоеваний и из добыч они посвящали на поддержание дома Господня.
1CHR|26|28|И все, что посвятил Самуил пророк, и Саул, сын Киса, и Авенир, сын Нира, и Иоав, сын Саруи, все посвященное [было] на руках у Шеломифа и братьев его.
1CHR|26|29|Из племени Ицгарова: Хенания и сыновья его [определены] на внешнее служение у Израильтян, писцами и судьями.
1CHR|26|30|Из племени Хевронова: Хашавия и братья его, люди мужественные, тысяча семьсот, имели надзор над Израилем по эту сторону Иордана к западу, по всяким делам [служения] Господня и по службе царской.
1CHR|26|31|У племени Хевронова Иерия [был] главою Хевронян, в их родах, в поколениях. В сороковой год царствования Давида они исчислены, и найдены между ними люди мужественные в Иазере Галаадском.
1CHR|26|32|И братья его, люди способные, две тысячи семьсот, были главы семейств. Их поставил царь Давид над коленом Рувимовым и Гадовым и полуколеном Манассииным, по всем делам Божиим и делам царя.
1CHR|27|1|Вот сыны Израилевы по числу их, главы семейств, тысяченачальники и стоначальники и управители, которые по отделениям служили царю во всех делах, приходя и отходя каждый месяц, во все месяцы года. В каждом отделении было их по двадцать четыре тысячи.
1CHR|27|2|Над первым отделением, для первого месяца, [начальствовал] Иашовам, сын Завдиила; в его отделении было двадцать четыре тысячи;
1CHR|27|3|он [был] из сынов Фареса, главный над всеми военачальниками в первый месяц.
1CHR|27|4|Над отделением второго месяца был Додай Ахохиянин; в отделении его был и князь Миклоф, и в его отделении было двадцать четыре тысячи.
1CHR|27|5|Третий главный военачальник, для третьего месяца, Ванея, сын Иодая, священника, и в его отделении было двадцать четыре тысячи:
1CHR|27|6|этот Ванея – [один] из тридцати храбрых и [начальник] над ними, и в его отделе [находился] Аммизавад, сын его.
1CHR|27|7|Четвертый, для четвертого месяца, был Асаил, брат Иоава, и по нем Завадия, сын его, и в его отделении двадцать четыре тысячи.
1CHR|27|8|Пятый, для пятого месяца, князь Шамгуф Израхитянин, и в его отделении двадцать четыре тысячи.
1CHR|27|9|Шестой, для шестого месяца, Ира, сын Иккеша, Фекоянин, и в его отделении двадцать четыре тысячи.
1CHR|27|10|Седьмой, для седьмого месяца, Хелец Пелонитянин, из сынов Ефремовых, и в его отделении двадцать четыре тысячи.
1CHR|27|11|Восьмой, для восьмого месяца, Совохай Хушатянин, из племени Зары, и в его отделении двадцать четыре тысячи.
1CHR|27|12|Девятый, для девятого месяца, Авиезер Анафофянин, из сыновей Вениаминовых, и в его отделении двадцать четыре тысячи.
1CHR|27|13|Десятый, для десятого месяца, Магарай Нетофафянин, из племени Зары, и в его отделении двадцать четыре тысячи.
1CHR|27|14|Одиннадцатый, для одиннадцатого месяца, Ванея Пирафонянин, из сынов Ефремовых, и в его отделении двадцать четыре тысячи.
1CHR|27|15|Двенадцатый, для двенадцатого месяца, Хелдай Нетофафянин, из потомков Гофониила, и в его отделении двадцать четыре тысячи.
1CHR|27|16|А над коленами Израилевыми, – у Рувимлян главным начальником [был] Елиезер, сын Зихри; у Симеона – Сафатия, сын Маахи;
1CHR|27|17|у Левия – Хашавия, сын Кемуила; у Аарона – Садок;
1CHR|27|18|у Иуды – Елиав, из братьев Давида; у Иссахара – Омри, сын Михаила;
1CHR|27|19|у Завулона – Ишмаия, сын Овадии; у Неффалима – Иеримоф, сын Азриила;
1CHR|27|20|у сыновей Ефремовых – Осия, сын Азазии; у полуколена Манассиина – Иоиль, сын Федаии;
1CHR|27|21|у полуколена Манассии в Галааде – Иддо, сын Захарии; у Вениамина – Иаасиил, сын Авенира;
1CHR|27|22|у Дана – Азариил, сын Иерохама. Вот вожди колен Израилевых.
1CHR|27|23|Давид не делал счисления тех, которые были от двадцати лет и ниже, потому что Господь сказал, что Он умножит Израиля, как звезды небесные.
1CHR|27|24|Иоав, сын Саруи, начал делать счисление, но не кончил. И был за это гнев Божий на Израиля, и не вошло то счисление в летопись царя Давида.
1CHR|27|25|Над сокровищами царскими был Азмавеф, сын Адиилов, а над запасами в поле, в городах, и в селах и в башнях – Ионафан, сын Уззии;
1CHR|27|26|над занимающимися полевыми работами, земледелием – Езрий, сын Хелува;
1CHR|27|27|над виноградниками – Шимей из Рамы, а над запасами вина в виноградниках – Завдий из Шефама;
1CHR|27|28|над маслинами и смоковницами в долине – Баал–Ханан Гедеритянин, а над запасами деревянного масла – Иоас;
1CHR|27|29|над крупным скотом, пасущимся в Шароне – Шитрай Шаронянин, а над скотом в долинах – Шафат, сын Адлая;
1CHR|27|30|над верблюдами – Овил Исмаильтянин; над ослицами – Иехдия Меронифянин;
1CHR|27|31|над мелким скотом – Иазиз Агаритянин. Все эти были начальниками над имением, которое [было] у царя Давида.
1CHR|27|32|Ионафан, дядя Давидов, [был] советником, человек умный и писец; Иехиил, сын Хахмониев, [был] при сыновьях царя;
1CHR|27|33|Ахитофел [был] советником царя; Хусий Архитянин – другом царя;
1CHR|27|34|после же Ахитофела Иодай, сын Ванеи, и Авиафар, а Иоав был военачальником у царя.
1CHR|28|1|И собрал Давид в Иерусалим всех вождей Израильских, начальников колен и начальников отделов, служивших царю, и тысяченачальников, и стоначальников, и заведывавших всем имением и стадами царя и сыновей его с евнухами, военачальников и всех храбрых мужей.
1CHR|28|2|И стал Давид царь на ноги свои и сказал: послушайте меня, братья мои и народ мой! [было] у меня на сердце построить дом покоя для ковчега завета Господня и в подножие ногам Бога нашего, и [потребное] для строения я приготовил.
1CHR|28|3|Но Бог сказал мне: не строй дома имени Моему, потому что ты человек воинственный и проливал кровь.
1CHR|28|4|Однакоже избрал Господь Бог Израилев меня из всего дома отца моего, чтоб быть [мне] царем над Израилем вечно, потому что Иуду избрал Он князем, а в доме Иуды дом отца моего, а из сыновей отца моего меня благоволил поставить царем над всем Израилем,
1CHR|28|5|из всех же сыновей моих, – ибо много сыновей дал мне Господь, – Он избрал Соломона, сына моего, сидеть на престоле царства Господня над Израилем,
1CHR|28|6|и сказал мне: Соломон, сын твой, построит дом Мой и дворы Мои, потому что Я избрал его Себе в сына, и Я буду ему Отцом;
1CHR|28|7|и утвержу царство его на веки, если он будет тверд в исполнении заповедей Моих и уставов Моих, как до сего дня.
1CHR|28|8|И теперь пред очами всего Израиля, собрания Господня, и во уши Бога нашего [говорю]: соблюдайте и держитесь всех заповедей Господа Бога вашего, чтобы владеть вам сею доброю землею и оставить ее после себя в наследство детям своим на век;
1CHR|28|9|и ты, Соломон, сын мой, знай Бога отца твоего и служи Ему от всего сердца и от всей души, ибо Господь испытует все сердца и знает все движения мыслей. Если будешь искать Его, то найдешь Его, а если оставишь Его, Он оставит тебя навсегда.
1CHR|28|10|Смотри же, когда Господь избрал тебя построить дом для святилища, будь тверд и делай.
1CHR|28|11|И отдал Давид Соломону, сыну своему, чертеж притвора и домов его, и кладовых его, и горниц его, и внутренних покоев его, и дома для ковчега,
1CHR|28|12|и чертеж всего, что было у него на душе, дворов дома Господня и всех комнат кругом, сокровищниц дома Божия и сокровищниц вещей посвященных,
1CHR|28|13|и священнических и левитских отделений, и всякого служебного дела в доме Господнем, и всех служебных сосудов дома Господня,
1CHR|28|14|золотых вещей, с [означением] веса, для всякого из служебных сосудов, всех вещей серебряных, с [означением] веса, для всякого из сосудов служебных.
1CHR|28|15|И дал золота для светильников и золотых лампад их, с означением веса каждого из светильников и лампад его, также светильников серебряных, с означением веса каждого из светильников и лампад его, смотря по служебному назначению каждого светильника;
1CHR|28|16|и золота для столов предложения хлебов, для каждого [золотого] стола, и серебра для столов серебряных,
1CHR|28|17|и вилок, и чаш и кропильниц из чистого золота, и золотых блюд, с означением веса каждого блюда, и серебряных блюд, с означением веса каждого блюда,
1CHR|28|18|и для жертвенника курения из литого золота с означением веса, и устройства колесницы с золотыми херувимами, распростирающими [крылья] и покрывающими ковчег завета Господня.
1CHR|28|19|Все сие в письмени от Господа, [говорил Давид, как] Он вразумил меня на все дела постройки.
1CHR|28|20|И сказал Давид сыну своему Соломону: будь тверд и мужествен, и приступай к делу, не бойся и не ужасайся, ибо Господь Бог, Бог мой, с тобою; Он не отступит от тебя и не оставит тебя, доколе не совершишь всего дела, требуемого для дома Господня.
1CHR|28|21|И вот отделы священников и левитов, для всякой службы при Доме Божием. И у тебя есть для всякого дела усердные люди, искусные для всякой работы, и начальники и весь народ [готовы] на все твои приказания.
1CHR|29|1|И сказал царь Давид всему собранию: Соломон, сын мой, которого одного избрал Бог, молод и малосилен, а дело сие велико, потому что не для человека здание сие, а для Господа Бога.
1CHR|29|2|Всеми силами я заготовил для дома Бога моего золото для золотых вещей и серебро для серебряных, и медь для медных, железо для железных, и дерева для деревянных, камни оникса и [камни] вставные, камни красивые и разноцветные, и всякие дорогие камни, и множество мрамора;
1CHR|29|3|и еще по любви моей к дому Бога моего, есть у меня сокровище собственное из золота и серебра, [и его] я отдаю для дома Бога моего, сверх всего, что заготовил я для святого дома:
1CHR|29|4|три тысячи талантов золота, золота Офирского, и семь тысяч талантов серебра чистого, для обложения стен в домах,
1CHR|29|5|для каждой из золотых вещей, и для каждой из серебряных, и для всякого изделия рук художнических. Не поусердствует ли [еще] кто жертвовать сегодня для Господа?
1CHR|29|6|И стали жертвовать начальники семейств и начальники колен Израилевых, и начальники тысяч и сотен, и начальники над имениями царя.
1CHR|29|7|И дали на устроение дома Божия пять тысяч талантов и десять тысяч драхм золота, и серебра десять тысяч талантов, и меди восемнадцать тысяч талантов, и железа сто тысяч талантов.
1CHR|29|8|И у кого нашлись [дорогие] камни, те отдавали и их в сокровищницу дома Господня, на руки Иехиилу Герсонитянину.
1CHR|29|9|И радовался народ усердию их, потому что они от всего сердца жертвовали Господу, также и царь Давид весьма радовался.
1CHR|29|10|И благословил Давид Господа пред всем собранием, и сказал Давид: благословен Ты, Господи Боже Израиля, отца нашего, от века и до века!
1CHR|29|11|Твое, Господи, величие, и могущество, и слава, и победа и великолепие, и все, [что] на небе и на земле, [Твое]: Твое, Господи, царство, и Ты превыше всего, как Владычествующий.
1CHR|29|12|И богатство и слава от лица Твоего, и Ты владычествуешь над всем, и в руке Твоей сила и могущество, и во власти Твоей возвеличить и укрепить все.
1CHR|29|13|И ныне, Боже наш, мы славословим Тебя и хвалим величественное имя Твое.
1CHR|29|14|Ибо кто я и кто народ мой, что мы имели возможность так жертвовать? Но от Тебя все, и от руки Твоей [полученное] мы отдали Тебе,
1CHR|29|15|потому что странники мы пред Тобою и пришельцы, как и все отцы наши, как тень дни наши на земле, и нет ничего прочного.
1CHR|29|16|Господи Боже наш! все это множество, которое приготовили мы для построения дома Тебе, святому имени Твоему, от руки Твоей оно, и все Твое.
1CHR|29|17|Знаю, Боже мой, что Ты испытуешь сердце и любишь чистосердечие; я от чистого сердца моего пожертвовал все сие, и ныне вижу, что и народ Твой, здесь находящийся, с радостью жертвует Тебе.
1CHR|29|18|Господи, Боже Авраама, Исаака и Израиля, отцов наших! сохрани сие навек, [сие] расположение мыслей сердца народа Твоего, и направь сердце их к Тебе.
1CHR|29|19|Соломону же, сыну моему, дай сердце правое, чтобы соблюдать заповеди Твои, откровения Твои и уставы Твои, и исполнить все это и построить здание, для которого я сделал приготовление.
1CHR|29|20|И сказал Давид всему собранию: благословите Господа Бога нашего. – И благословило все собрание Господа Бога отцов своих, и пало, и поклонилось Господу и царю.
1CHR|29|21|И принесли Господу жертвы, и вознесли всесожжения Господу, на другой после сего день: тысячу тельцов, тысячу овнов, тысячу агнцев с их возлияниями, и множество жертв от всего Израиля.
1CHR|29|22|И ели и пили пред Господом в тот день, с великою радостью; и в другой раз воцарили Соломона, сына Давидова, и помазали пред Господом в правителя верховного, а Садока во священника.
1CHR|29|23|И сел Соломон на престоле Господнем, как царь, вместо Давида, отца своего, и был благоуспешен, и весь Израиль повиновался ему.
1CHR|29|24|И все начальники и сильные, также и все сыновья царя Давида подчинились Соломону царю.
1CHR|29|25|И возвеличил Господь Соломона пред очами всего Израиля, и даровал ему славу царства, какой не имел прежде его ни один царь у Израиля.
1CHR|29|26|И Давид, сын Иессеев, царствовал над всем Израилем.
1CHR|29|27|Времени царствования его над Израилем [было] сорок лет: в Хевроне царствовал он семь лет, и в Иерусалиме царствовал тридцать три [года].
1CHR|29|28|И умер в доброй старости, насыщенный жизнью, богатством и славою; и воцарился Соломон, сын его, вместо него.
1CHR|29|29|Дела царя Давида, первые и последние, описаны в записях Самуила провидца и в записях Нафана пророка и в записях Гада прозорливца,
1CHR|29|30|равно и все царствование его, и мужество его, и происшествия, случившиеся с ним и с Израилем и со всеми земными царствами.
