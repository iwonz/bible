NEH|1|1|Verba Nehemiae filii Hacha liae. Et factum est in mense Ca sleu, anno vicesimo, et ego eram in castro Susan.
NEH|1|2|Et venit Hanani unus de fratribus meis, ipse et viri ex Iuda; et interrogavi eos de Iudaeis, qui salvati erant et supererant de captivitate, et de Ierusalem.
NEH|1|3|Et dixerunt mihi: " Superstites, qui supererant de captivitate ibi in provincia, in afflictione magna sunt et in opprobrio; et murus Ierusalem dissipatus est, et portae eius combustae sunt igne ".
NEH|1|4|Cumque audissem verba huiuscemodi, sedi et flevi et luxi diebus multis; ieiunabam et orabam ante faciem Dei caeli.
NEH|1|5|Et dixi: " Quaeso, Domine, Deus caeli, Deus fortis, magne atque terribilis, qui custodis pactum et misericordiam cum his, qui te diligunt et custodiunt mandata tua;
NEH|1|6|fiat auris tua auscultans, et oculi tui aperti, ut audias orationem servi tui, quam ego oro coram te hodie, die et nocte pro filiis Israel servis tuis, et confiteor pro peccatis filiorum Israel, quibus peccaverunt tibi. Ego quoque et domus patris mei peccavimus,
NEH|1|7|delinquentes deliquimus contra te et non custodivimus praecepta et mandata et iudicia, quae praecepisti Moysi famulo tuo.
NEH|1|8|Memento verbi, quod mandasti Moysi servo tuo dicens: "Cum transgressi fueritis, ego dispergam vos in populos;
NEH|1|9|si autem revertamini ad me et custodiatis praecepta mea et faciatis ea, etiamsi abducti fueritis in extrema caeli, inde congregabo vos et reducam in locum quem elegi, ut habitaret nomen meum ibi".
NEH|1|10|Ipsi enim sunt servi tui et populus tuus, quos redemisti in fortitudine tua magna et in manu tua valida.
NEH|1|11|Obsecro, Domine, sit auris tua attendens ad orationem servi tui et ad orationem servorum tuorum, qui volunt timere nomen tuum; et fac servum tuum prosperari hodie et da ei gratiam ante virum hunc ". Ego enim eram pincerna regis.
NEH|2|1|Factum est autem in mense Nisan, anno vicesimo Artaxerxis regis, dum biberet, levavi vinum et dedi regi; non enim eram ingratus coram eo.
NEH|2|2|Dixitque mihi rex: " Quare vultus tuus tristis est, cum te aegrotum non videam? Nihil est aliud nisi tristitia cordis ". Et timui valde
NEH|2|3|et dixi regi: " Rex, in aeternum vive! Quare non maereat vultus meus, quia civitas sepulcrorum patrum meorum deserta est, et portae eius combustae sunt igne? ".
NEH|2|4|Et ait mihi rex: " Pro qua re postulas? ". Et oravi Deum caeli
NEH|2|5|et dixi ad regem: " Si videtur regi bonum, et si placet servus tuus ante faciem tuam, ut mittas me in Iudaeam ad civitatem sepulcrorum patrum meorum, et aedificabo eam ".
NEH|2|6|Dixitque mihi rex, et regina sedebat iuxta eum: " Usque ad quod tempus erit iter tuum, et quando reverteris? ". Et placuit regi mittere me; et constitui ei tempus.
NEH|2|7|Et dixi regi: " Si regi videtur bonum, epistulae dentur mihi ad duces regionis trans flumen, ut me transire permittant, donec veniam in Iudaeam;
NEH|2|8|et epistulam ad Asaph custodem saltus regis, ut det mihi ligna, ut contignare possim portas turris domus et muri civitatis et domus, in qua habitabo ". Et dedit mihi rex, quia manus Dei mei bona super me.
NEH|2|9|Et veni ad duces regionis trans flumen dedique eis epistulas regis. Miserat autem rex mecum principes militum et equites.
NEH|2|10|Et audierunt Sanaballat Horonites et Thobias servus Ammanites et contristati sunt afflictione magna, quod venisset homo, qui quaereret prosperitatem filiorum Israel.
NEH|2|11|Et veni Ierusalem et eram ibi tribus diebus.
NEH|2|12|Et surrexi nocte ego, et viri pauci mecum, et non indicavi cuiquam quid Deus meus dedisset in corde meo, ut facerem in Ierusalem; et iumentum non erat mecum, nisi animal cui sedebam.
NEH|2|13|Et egressus sum per portam Vallis nocte et ad fontem Draconis et portam Sterquilinii et considerabam murum Ierusalem dissipatum et portas eius consumptas igne.
NEH|2|14|Et transivi ad portam Fontis et ad piscinam Regis, et non erat locus iumento cui sedebam, ut transiret.
NEH|2|15|Et ascendi per torrentem nocte et considerabam murum; et iterum veni ad portam Vallis et reversus sum.
NEH|2|16|Magistratus autem nesciebant quo abissem aut quid ego facerem, sed et Iudaeis et sacerdotibus et optimatibus et magistratibus et reliquis, qui faciebant opus, usque ad id loci nihil indicaveram.
NEH|2|17|Et dixi eis: " Vos nostis afflictionem, in qua sumus, quia Ierusalem deserta est, et portae eius consumptae sunt igne; venite et aedificemus murum Ierusalem et non simus ultra opprobrium ".
NEH|2|18|Et indicavi eis quod manus Dei mei bona esset super me et verba regis, quae locutus esset mihi, et dixerunt: " Surgamus et aedificemus! ". Et confortatae sunt manus eorum in bonum.
NEH|2|19|Audierunt autem Sanaballat Horonites et Thobias servus Ammanites et Gosem Arabs et subsannaverunt nos et despexerunt dixeruntque: " Quae est haec res, quam facitis? Numquid contra regem vos rebellatis? ".
NEH|2|20|Et dedi eis responsum dicens: " Deus caeli ipse nos facit prosperari, et nos servi eius sumus; surgamus et aedificemus. Vobis autem non est pars et ius et memoria in Ierusalem ".
NEH|3|1|Et surrexit Eliasib sacerdos magnus et fratres eius sacerdotes et aedificaverunt portam Gregis; contignaverunt eam et statuerunt valvas eius et usque ad turrim Meah et turrim Hananeel.
NEH|3|2|Et iuxta eos aedificaverunt viri Iericho, et iuxta eos aedificavit Zacchur filius Imri.
NEH|3|3|Portam autem Piscium aedificaverunt filii Asnaa; ipsi contignaverunt eam et statuerunt valvas eius et seras et vectes.
NEH|3|4|Et iuxta eos restauravit Meremoth filius Uriae filii Accos, et iuxta eum restauravit Mosollam filius Barachiae filii Mesezabel, et iuxta eum restauravit Sadoc filius Baana,
NEH|3|5|et iuxta eum restauraverunt Thecueni; optimates autem eorum non supposuerunt colla sua in opere Domini sui.
NEH|3|6|Et portam Veterem restauraverunt Ioiada filius Phasea et Mosollam filius Besodia; ipsi contignaverunt eam et statuerunt valvas eius et seras et vectes.
NEH|3|7|Et iuxta eos restauraverunt Meltias Gabaonites et Iadon Meronathites, viri de Gabaon et Maspha, qui erant ad solium ducis, qui erat in regione trans flumen;
NEH|3|8|et iuxta eos restauravit Oziel filius Araia de aurificibus, et iuxta eum restauravit Hananias de pigmentariis et firmaverunt Ierusalem usque ad murum latiorem.
NEH|3|9|Et iuxta eum restauravit Raphaia filius Hur, princeps dimidiae partis vici Ierusalem;
NEH|3|10|et iuxta eum restauravit Iedaia filius Haromaph contra domum suam, et iuxta eum restauravit Hattus filius Hasabneia.
NEH|3|11|Alteram partem restauravit Melchias filius Harim et Hassub filius Phahathmoab usque ad turrim Furnorum.
NEH|3|12|Et iuxta eos restauravit Sellum filius Alohes, princeps mediae partis vici Ierusalem, ipse et filiae eius.
NEH|3|13|Portam Vallis restauravit Hanun et habitatores Zanoa; ipsi aedificaverunt eam et statuerunt valvas eius et seras et vectes et mille cubitos in muro usque ad portam Sterquilinii.
NEH|3|14|Et portam Sterquilinii restauravit Melchias filius Rechab, princeps vici Bethcharem; ipse aedificavit eam et statuit valvas eius et seras et vectes.
NEH|3|15|Et portam Fontis restauravit Sellum filius Cholhoza princeps pagi Maspha; ipse aedificavit eam et texit et statuit valvas eius et seras et vectes et murum piscinae Siloae iuxta hortum regis et usque ad gradus, qui descendunt de civitate David.
NEH|3|16|Post eum restauravit Nehemias filius Azboc princeps dimidiae partis vici Bethsur usque contra sepulcra David et usque ad piscinam, quae repleta est, et usque ad domum Fortium.
NEH|3|17|Post eum restauraverunt Levitae, Rehum filius Bani; iuxta eum restauravit Hasabias princeps dimidiae partis vici Ceilae pro vico suo;
NEH|3|18|post eum aedificaverunt fratres eorum Bavai filius Henadad princeps dimidiae partis vici Ceilae.
NEH|3|19|Et restauravit iuxta eum Ezer filius Iesua princeps Maspha mensuram alteram contra ascensum armentarii in angulo.
NEH|3|20|Post eum restauravit Baruch filius Zachai mensuram alteram ab angulo usque ad portam domus Eliasib sacerdotis magni.
NEH|3|21|Post eum restauravit Meremoth filius Uriae filii Aecos mensuram secundam a porta domus Eliasib usque ad extremitatem domus Eliasib.
NEH|3|22|Et post eum restauraverunt sacerdotes viri de campestribus.
NEH|3|23|Post eos restauravit Beniamin et Hassub contra domum suam; post eos restauravit Azarias filius Maasiae filii Ananiae iuxta domum suam.
NEH|3|24|Post eum restauravit Bennui filius Henadad mensuram alteram a domo Azariae usque ad angulum et flexuram.
NEH|3|25|Phalel filius Ozi contra angulum turris, quae eminet de domo regis excelsa in atrio carceris; post eum Phadaia filius Pharos restauravit
NEH|3|26|usque contra portam Aquarum ad orientem et turrim, quae prominebat.
NEH|3|27|Post eum restauraverunt Thecueni mensuram alteram a regione contra magnam turrim eminentem usque ad murum templi.
NEH|3|28|Sursum autem a porta Equorum restauraverunt sacerdotes, unusquisque contra domum suam.
NEH|3|29|Post eos restauravit Sadoc filius Emmer contra domum suam; et post eum restauravit Semeia filius Secheniae custos portae orientalis.
NEH|3|30|Post eum restauravit Hanania filius Selemiae et Hanun filius Seleph sextus mensuram alteram. Post eum restauravit Mosollam filius Barachiae contra cellam suam.
NEH|3|31|Post eum restauravit Melchias de aurificibus usque ad domum oblatorum et mercatorum, contra portam Iudicialem, et usque ad cenaculum anguli;
NEH|3|32|et inter cenaculum anguli et portam Gregis restauraverunt aurifices et negotiatores.
NEH|3|33|Factum est autem, cum audisset Sanaballat quod aedificaremus murum, iratus est et indignatus est nimis et subsannavit Iudaeos
NEH|3|34|et dixit coram fratribus suis et optimatibus Samariae: " Quid Iudaei faciunt imbecilles? Num hoc conceditur eis? Num, quia sacrificant, complebunt in una die? Numquid vivificare poterunt lapides de acervis pulveris, qui combusti sunt? ".
NEH|3|35|Sed et Thobias Ammanites, qui erat ad latus eius, ait: " Sine aedificare; si ascenderit vulpes, diruet murum eorum lapideum ".
NEH|3|36|Audi, Deus noster, quia facti sumus irrisio! Converte contumeliam eorum super caput eorum et da eos in irrisionem in terra captivitatis!
NEH|3|37|Ne operias iniquitatem eorum, et peccatum eorum coram facie tua non deleatur, quia offenderunt te coram aedificantibus.
NEH|3|38|Itaque aedificavimus murum, et compositus est totus murus usque ad partem dimidiam, et populus dabat cor suum, ut operaretur.
NEH|4|1|Factum est autem cum audisset Sanaballat et Thobias et Arabes et Ammanitae et Azotii quod prosperaretur restauratio muri Ierusalem et quod coepissent interrupta concludi, irati sunt nimis;
NEH|4|2|et conspiraverunt omnes pariter, ut venirent et pugnarent contra Ierusalem et facerent confusionem.
NEH|4|3|Et oravimus Deum nostrum et posuimus custodiam die ac nocte contra eos.
NEH|4|4|Dixit autem Iudas: " Debilitata est fortitudo portantis, et humus nimia est; et nos non poterimus aedificare murum ".
NEH|4|5|Et dixerunt hostes nostri: " Nesciant et ignorent, donec veniamus in medium eorum et interficiamus eos et cessare faciamus opus ".
NEH|4|6|Factum est autem venientibus Iudaeis, qui habitabant iuxta eos, et dicentibus nobis per decem vices ex omnibus locis, quibus venerant ad nos,
NEH|4|7|statuimus nos in inferioribus post murum in locis apertis, et ordinavi populum secundum familias cum gladiis suis et lanceis suis et arcubus suis.
NEH|4|8|Et perspexi atque surrexi, et aio ad optimates et magistratus et ad reliquam partem vulgi: " Nolite timere a facie eorum; Domini magni et terribilis mementote et pugnate pro fratribus vestris, filiis vestris et filiabus vestris et uxoribus vestris et domibus vestris ".
NEH|4|9|Factum est autem cum audissent inimici nostri nuntiatum esse nobis, dissipavit Deus consilium eorum, et reversi sumus omnes ad murum, unusquisque ad opus suum.
NEH|4|10|Et factum est a die illa, media pars iuvenum meorum faciebat opus, et media tenebat lanceas et scuta et arcus et loricas, et principes post omnem domum Iudae.
NEH|4|11|Aedificantium in muro et portantium onera et imponentium, una manu sua faciebat opus et altera tenebat gladium;
NEH|4|12|aedificantium enim unusquisque gladio erat accinctus renes, et sic aedificabant; et, qui clangebat bucina, iuxta me.
NEH|4|13|Et dixi ad optimates et ad magistratus et ad reliquam partem vulgi: " Opus grande est et latum, et nos separati sumus in muro procul alter ab altero;
NEH|4|14|in loco quocumque audieritis clangorem tubae, illuc concurrite ad nos. Deus noster pugnabit pro nobis ".
NEH|4|15|Et sic nos fecimus opus, et media pars nostrum tenebat lanceas ab ascensu aurorae, donec egrediantur astra.
NEH|4|16|In tempore quoque illo dixi populo: " Unusquisque cum puero suo pernoctet in medio Ierusalem; et erit nobis custodia per noctem, et opus per diem ".
NEH|4|17|Ego autem et fratres mei et pueri mei et custodes, qui erant post me, non deponebamus vestimenta nostra; unusquisque tenebat gladium in dextera sua.
NEH|5|1|Et factus est clamor populi et uxorum eius magnus adversus fratres suos Iudaeos.
NEH|5|2|Et erant qui dicerent: " Filios nostros et filias nostras pignoravimus, ut acciperemus frumentum et comederemus et viveremus! ".
NEH|5|3|Et erant qui dicerent: " Agros nostros et vineas et domos nostras opposuimus, ut acciperemus frumentum in fame! ".
NEH|5|4|Et alii dicebant: " Mutuo sumpsimus pecunias in tributa regis pro agris nostris et vineis nostris.
NEH|5|5|Et nunc sicut caro fratrum nostrorum sic caro nostra est, et sicut filii eorum ita et filii nostri; ecce nos subiugamus filios nostros et filias nostras in servitutem, et de filiabus nostris quaedam iam in servitute subiugatae sunt, nec habemus unde possint redimi, quia agros nostros et vineas nostras alii possident ".
NEH|5|6|Et iratus sum nimis, cum audissem clamorem eorum secundum verba haec.
NEH|5|7|Cogitavique in corde meo et increpavi optimates et magistratus et dixi eis: " Usuras singuli a fratribus vestris exigitis! ". Et congregavi adversum eos contionem magnam
NEH|5|8|et dixi eis: " Nos, ut scitis, redemimus fratres nostros Iudaeos, qui venditi fuerant gentibus, secundum possibilitatem nostram; quin potius et vos vendetis fratres vestros, ut vendentur nobis? ". Et siluerunt nec invenerunt quid responderent.
NEH|5|9|Dixique ad eos: " Non est bona res, quam facitis. Quare non in timore Dei nostri ambulatis, ne exprobretur nobis a gentibus inimicis nostris?
NEH|5|10|Et ego et fratres mei et pueri mei commodavimus plurimis pecuniam et frumentum; non repetamus usuras istas.
NEH|5|11|Reddite eis hodie agros suos et vineas suas et oliveta sua et domos suas et centesimam pecuniae frumenti vini et olei, quam exigere soletis ab eis ".
NEH|5|12|Et dixerunt: " Reddemus et ab eis nihil quaeremus; sicque faciemus, ut loqueris ". Et vocavi sacerdotes et feci eos iurare, ut facerent, sicut dictum erat.
NEH|5|13|Insuper excussi sinum meum et dixi: " Sic excutiat Deus omnem virum, qui non compleverit verbum istud, de domo sua et de laboribus suis; sic excutiatur et vacuus fiat! ". Et dixit universa multitudo: " Amen! ". Et laudaverunt Deum. Fecit ergo populus, sicut erat dictum.
NEH|5|14|A die autem illa, qua praeceperat rex mihi, ut essem dux in terra Iudae, ab anno vicesimo usque ad annum tricesimum secundum Artaxerxis regis, per annos duodecim ego et fratres mei annonas, quae ducibus debebantur, non comedimus.
NEH|5|15|Duces autem priores, qui fuerant ante me, gravaverunt populum et acceperunt ab eis cotidie pro pane siclos argenti quadraginta; sed et ministri eorum depresserunt populum. Ego autem non feci ita propter timorem Dei,
NEH|5|16|quin potius in opere muri restauravi et agrum non emi; et omnes pueri mei congregati ad opus erant.
NEH|5|17|Iudaei quoque et magistratus, centum quinquaginta viri, et qui veniebant ad nos de gentibus, quae in circuitu nostro sunt, in mensa mea erant.
NEH|5|18|Parabatur autem mihi per dies singulos bos unus, arietes sex electi, exceptis volatilibus; et inter dies decem vina diversa multa. Insuper et annonas ducatus mei non quaesivi; gravis enim erat servitus populi huius.
NEH|5|19|Memento mei, Deus meus, in bonum, secundum omnia, quae feci populo huic.
NEH|6|1|Factum est autem cum audisset Sanaballat et Thobias et Gosem Arabs et ceteri inimici nostri, quod aedificassem ego murum, et non esset in ipso residua interruptio - usque ad tempus autem illud valvas non posueram in portis -
NEH|6|2|miserunt Sanaballat et Gosem ad me dicentes: " Veni, et conveniamus in Cephirim in campo Ono ". Ipsi autem cogitabant, ut facerent mihi malum.
NEH|6|3|Misi ergo ad eos nuntios dicens: " Opus grande ego facio et non possum descendere; cur cessare oportet opus, si desistero et descendero ad vos?.
NEH|6|4|Miserunt autem ad me secundum verbum hoc per quattuor vices, et respondi eis iuxta sermonem priorem.
NEH|6|5|Et misit ad me Sanaballat iuxta verbum prius quinta vice puerum suum, et epistulam non obsignatam habebat in manu sua, in qua erat scriptum:
NEH|6|6|" In gentibus auditum est, et Gosem dixit quod tu et Iudaei cogitetis rebellare, et propterea aedifices murum et levare te velis super eos regem; iuxta hanc vocem
NEH|6|7|et prophetas posueris, qui praedicent de te in Ierusalem dicentes: "Rex in Iudaea est!". Nunc autem auditurus est rex verba haec; idcirco nunc veni, ut ineamus consilium pariter ".
NEH|6|8|Et misi ad eum dicens: " Non est factum secundum verba haec, quae tu loqueris; de corde enim tuo tu componis haec ".
NEH|6|9|Omnes enim hi terrebant nos cogitantes: " Fatigabuntur manus eorum ab opere, et non complebitur ". Quam ob causam magis confortavi manus meas.
NEH|6|10|Et ingressus sum domum Semeiae filii Dalaiae filii Meetabel, ubi erat detentus. Qui ait: " Tractemus nobiscum in domo Dei, in medio templi, et claudamus portas aedis, quia venturi sunt, ut interficiant te; utique nocte venturi sunt ad occidendum te".
NEH|6|11|Et dixi: " Num quisquam similis mei fugit? Et quis ut ego ingredietur templum et vivet? Non ingrediar ".
NEH|6|12|Et intellexi quod Deus non misisset eum, sed quasi vaticinans locutus esset ad me, quia Thobias et Sanaballat conduxerant eum.
NEH|6|13|Acceperat enim pretium, ut territus sic agerem et peccarem, et haberent malum, quod exprobrarent mihi.
NEH|6|14|Memento, Deus meus, Thobiae et Sanaballat iuxta opera eorum talia, sed et Noadiae prophetae et ceterorum prophetarum, qui terrebant me!
NEH|6|15|Completus est autem murus vicesimo quinto die mensis Elul, quinquaginta duobus diebus.
NEH|6|16|Factum est ergo, cum audissent omnes inimici nostri, et vidissent universae gentes, quae erant in circuitu nostro, ut conciderent intra semetipsos et scirent quod a Deo factum esset opus hoc.
NEH|6|17|Sed et in diebus illis, multae optimatum Iudaeorum epistulae mittebantur ad Thobiam, et a Thobia veniebant ad eos.
NEH|6|18|Multi enim in Iudaea coniurationem fecerunt cum eo, quia gener erat Secheniae filii Area, et Iohanan filius eius acceperat filiam Mosollam filii Barachiae.
NEH|6|19|Sed et laudabant eum coram me et verba mea nuntiabant ei; et Thobias mittebat epistulas, ut terreret me.
NEH|7|1|Postquam autem aedificatus est murus, et posui valvas et recen sui ianitores et cantores et Levitas,
NEH|7|2|praeposui Hanani fratrem meum et Hananiam principem arcis supra Ierusalem - ipse enim quasi vir verax et timens Deum plus ceteris videbatur -
NEH|7|3|et dixi eis: " Non aperiantur portae Ierusalem usque ad calorem solis. Dum adhuc calor permanet, claudantur portae et oppilentur; et ponant custodes de habitatoribus Ierusalem, singulos per vices suas et unumquemque contra domum suam ".
NEH|7|4|Civitas autem erat lata nimis et grandis, et populus parvus in medio eius, et non erant domus aedificatae.
NEH|7|5|Deus autem meus dedit in corde meo, et congregavi optimates et magistratus et vulgus, ut recenserem eos; et inveni librum census eorum, qui ascenderant primum, et inventum est scriptum in eo:
NEH|7|6|Isti filii provinciae, qui ascenderunt de captivitate migrantium, quos transtulerat Nabuchodonosor rex Babylonis, et reversi sunt in Ierusalem et in Iudaeam unusquisque in civitatem suam.
NEH|7|7|Qui venerunt cum Zorobabel, Iesua, Nehemias, Azarias, Raamias, Nahamani, Mardochaeus, Belsan, Mespharath, Beguai, Nahum, Baana.Numerus virorum populi Israel:
NEH|7|8|filii Pharos duo milia centum septuaginta duo;
NEH|7|9|filii Saphatia trecenti septuaginta duo;
NEH|7|10|filii Area sescenti quinquaginta duo;
NEH|7|11|filii Phahathmoab, hi sunt filii Iesua et Ioab, duo milia octingenti decem et octo;
NEH|7|12|filii Elam mille ducenti quinquaginta quattuor;
NEH|7|13|filii Zethua octingenti quadraginta quinque;
NEH|7|14|filii Zachai septingenti sexaginta;
NEH|7|15|filii Bennui sescenti quadraginta octo;
NEH|7|16|filii Bebai sescenti viginti octo;
NEH|7|17|filii Azgad duo milia trecenti viginti duo;
NEH|7|18|filii Adonicam sescenti sexaginta septem;
NEH|7|19|filii Beguai duo milia sexaginta septem;
NEH|7|20|filii Adin sescenti quinquaginta quinque;
NEH|7|21|filii Ater, qui erant ex Ezechia, nonaginta octo;
NEH|7|22|filii Hasum trecenti viginti octo;
NEH|7|23|filii Besai trecenti viginti quattuor;
NEH|7|24|filii Hareph centum duodecim;
NEH|7|25|filii Gabaon nonaginta quinque;
NEH|7|26|filii Bethlehem et Netopha centum octoginta octo;
NEH|7|27|viri Anathoth centum viginti octo;
NEH|7|28|viri Bethazmaveth quadraginta duo;
NEH|7|29|viri Cariathiarim, Cephira et Beroth septingenti quadraginta tres;
NEH|7|30|viri Rama et Gabaa sescenti viginti unus;
NEH|7|31|viri Machmas centum viginti duo;
NEH|7|32|viri Bethel et Hai centum viginti tres;
NEH|7|33|viri Nabo alterius quinquaginta duo;
NEH|7|34|viri Elam alterius mille ducenti quinquaginta quattuor;
NEH|7|35|filii Harim trecenti viginti;
NEH|7|36|filii Iericho trecenti quadraginta quinque;
NEH|7|37|filii Lod, Hadid et Ono septingenti viginti unus;
NEH|7|38|filii Senaa tria milia nongenti triginta.
NEH|7|39|Sacerdotes: filii Iedaia de domo Iesua nongenti septuaginta tres;
NEH|7|40|filii Emmer mille quinquaginta duo;
NEH|7|41|filii Phassur mille ducenti quadraginta septem;
NEH|7|42|filii Harim mille decem et septem.
NEH|7|43|Levitae: filii Iesua, hi sunt filii Cadmihel, Bennui et Odoviae, septuaginta quattuor.
NEH|7|44|Cantores: filii Asaph centum quadraginta octo.
NEH|7|45|Ianitores: filii Sellum, filii Ater, filii Telmon, filii Accub, filii Hatita, filii Sobai, centum triginta octo.
NEH|7|46|Oblati: filii Siha, filii Hasupha, filii Tabbaoth,
NEH|7|47|filii Ceros, filii Siaa, filii Phadon,
NEH|7|48|filii Lebana, filii Hagaba, filii Selmai,
NEH|7|49|filii Hanan, filii Giddel, filii Gaher,
NEH|7|50|filii Raaia, filii Rasin, filii Necoda,
NEH|7|51|filii Gazam, filii Oza, filii Phasea,
NEH|7|52|filii Besai, filii Meunitarum, filii Nephusorum,
NEH|7|53|filii Bacbuc, filii Hacupha, filii Harhur,
NEH|7|54|filii Basluth, filii Mahida, filii Harsa,
NEH|7|55|filii Bercos, filii Sisara, filii Thema,
NEH|7|56|filii Nasia, filii Hatipha.
NEH|7|57|Filii servorum Salomonis: filii Sotai, filii Sophereth, filii Pheruda,
NEH|7|58|filii Iaala, filii Darcon, filii Giddel,
NEH|7|59|filii Saphatia, filii Hatil, filii Phochereth Hassebaim, filii Amon.
NEH|7|60|Omnes oblati et filii servorum Salomonis trecenti nonaginta duo.
NEH|7|61|Hi sunt autem, qui ascenderunt de Thelmela, Thelharsa, Cherub, Addon et Emmer et non potuerunt indicare domum patrum suorum et semen suum, utrum ex Israel essent:
NEH|7|62|filii Dalaia, filii Thobia, filii Necoda sescenti quadraginta duo.
NEH|7|63|Et de sacerdotibus: filii Hobia, filii Accos, filii Berzellai, qui accepit de filiabus Berzellai Galaaditis uxorem et vocatus est nomine eorum.
NEH|7|64|Hi quaesierunt tabulas genealogiae suae et non invenerunt; et eiecti sunt de sacerdotio;
NEH|7|65|dixitque praepositus eis, ut non manducarent de sanctificatis sanctuarii, donec staret sacerdos pro Urim et Tummim.
NEH|7|66|Omnis multitudo simul quadraginta duo milia trecenti sexaginta,
NEH|7|67|absque servis et ancillis eorum, qui erant septem milia trecenti triginta septem; insuper et cantores et cantatrices ducenti quadraginta quinque.
NEH|7|68|Equi eorum septingenti triginta sex, muli eorum ducenti quadraginta quinque,
NEH|7|69|cameli eorum quadringenti triginta quinque, asini sex milia septingenti viginti.
NEH|7|70|Nonnulli autem de principibus familiarum dederunt in opus: praepositus dedit in thesaurum auri drachmas mille, phialas quinquaginta, tunicas sacerdotales quingentas triginta;
NEH|7|71|et de principibus familiarum dederunt in thesaurum operis auri drachmas viginti milia et argenti minas duo milia ducentas.
NEH|7|72|Et quod dedit reliquus populus, auri drachmas viginti milia et argenti minas duo milia et tunicas sacerdotales sexaginta septem. Habitaverunt autem ibi sacerdotes et Levitae; ianitores autem et cantores et quidam de populo et oblati et omnis Israel habitaverunt in civitatibus suis.Et venerat mensis septimus; filii autem Israel erant in civitatibus suis.
NEH|8|1|Congregatusque est omnis populus quasi vir unus ad plateam, quae est ante portam Aquarum, et dixerunt Esdrae scribae, ut afferret librum legis Moysi, quam praece perat Dominus Israeli.
NEH|8|2|Attulit ergo Esdras sacerdos legem coram multitudine virorum et mulierum cunctisque, qui poterant intellegere, in die prima mensis septimi.
NEH|8|3|Et legit in eo in platea, quae erat ante portam Aquarum, de mane usque ad mediam diem in conspectu virorum et mulierum et eorum, qui intellegere poterant; et aures omnis populi erant erectae ad librum legis.
NEH|8|4|Stetit autem Esdras scriba super gradum ligneum, quem ad hoc fecerant; et steterunt iuxta eum Matthathias et Sema et Anaia et Uria et Helcia et Maasia ad dexteram eius, et ad sinistram Phadaia, Misael et Melchia et Hasum et Hasbadana, Zacharia et Mosollam.
NEH|8|5|Et aperuit Esdras librum coram omni populo - super universum quippe populum eminebat - et, cum aperuisset eum, stetit omnis populus.
NEH|8|6|Et benedixit Esdras Domino, Deo magno; et respondit omnis populus: " Amen, amen ", elevans manus suas. Et incurvati sunt et adoraverunt Deum proni in terram.
NEH|8|7|Porro Iesua et Bani et Serebia, Iamin, Accub, Sabethai, Hodia, Maasia, Celita, Azarias, Iozabad, Hanan, Phalaia et Levitae erudiebant populum in lege; populus autem stabat in gradu suo.
NEH|8|8|Et legerunt in libro legis Dei distincte et aperierunt sensum et explicaverunt lectionem.
NEH|8|9|Dixit autem Nehemias, ipse est praepositus, et Esdras sacerdos et scriba et Levitae instruentes populum universo populo: " Dies iste sanctificatus est Domino Deo nostro! Nolite lugere et nolite flere ". Flebat enim omnis populus, cum audiret verba legis.
NEH|8|10|Et dixit eis: " Ite, comedite pinguia et bibite mulsum et mittite partes his, qui non praeparaverunt sibi, quia sanctus dies Domini nostri est; et nolite contristari, gaudium etenim Domini est fortitudo vestra ".
NEH|8|11|Levitae autem silentium faciebant in omni populo dicentes: " Tacete, quia dies sanctus est, et nolite dolere ".
NEH|8|12|Abiit itaque omnis populus, ut comederet et biberet et mitteret partes et faceret laetitiam magnam, quia intellexerant verba, quae docuerat eos.
NEH|8|13|Et in die secundo congregati sunt principes familiarum universi populi, sacerdotes et Levitae ad Esdram scribam, ut intellegerent verba legis.
NEH|8|14|Et invenerunt scriptum in lege, quam praecepit Dominus per Moysen, ut habitent filii Israel in tabernaculis in die sollemni mense septimo
NEH|8|15|et ut praedicent et divulgent vocem in universis urbibus suis et in Ierusalem dicentes: " Egredimini in montem et afferte frondes olivae et frondes oleastri, frondes myrti et ramos palmarum et frondes ligni nemorosi, ut fiant tabernacula, sicut scriptum est ".
NEH|8|16|Et egressus est populus, et attulerunt feceruntque sibi tabernacula, unusquisque in domate suo et in atriis suis et in atriis domus Dei et in platea portae Aquarum et in platea portae Ephraim.
NEH|8|17|Fecit ergo universa ecclesia eorum, qui redierant de captivitate, tabernacula et habitaverunt in tabernaculis. Non enim fecerant a diebus Iosue filii Nun taliter filii Israel usque ad diem illum; et fuit laetitia magna nimis.
NEH|8|18|Legit autem in libro legis Dei per dies singulos, a die primo usque ad diem novissimum; et fecerunt sollemnitatem septem diebus et in die octavo conventum iuxta ordinationem.
NEH|9|1|In die autem vicesimo quarto mensis huius convenerunt filii Is rael in ieiunio et in saccis, et humus super eos.
NEH|9|2|Et separatum est semen filiorum Israel ab omni alienigena; et steterunt et confitebantur peccata sua et iniquitates patrum suorum.
NEH|9|3|Et consurrexerunt ad standum et legerunt in volumine legis Domini Dei sui per quartam partem diei; et per quartam partem confitebantur et adorabant Dominum Deum suum.
NEH|9|4|Surrexerunt autem super gradum Levitarum Iesua et Bani et Cadmihel, Sebania, Bunni, Serebia, Bani et Chanani et clamaverunt voce magna ad Dominum Deum suum.
NEH|9|5|Et dixerunt Levitae Iesua et Cadmihel, Bani, Hasabneia, Serebia, Hodia, Sebania, Phethahia: Surgite, benedicite Domino Deo vestroab aetemo usque in aeternum,et benedicant nomini gloriae tuae excelsosuper omnem benedictionem et laudem.
NEH|9|6|Tu ipse, Domine, solus;tu fecisti caelum et caelum caelorumet omnem exercitum eorum,terram et universa, quae in ea sunt, maria et omnia, quae in eis sunt;et tu vivificas omnia haec,et exercitus caeli te adorat.
NEH|9|7|Tu ipse, Domine Deus, qui elegisti Abramet eduxisti eum de Ur Chaldaeorumet posuisti nomen eius Abraham.
NEH|9|8|Et invenisti cor eius fidele coram teet percussisti cum eo foedus,ut dares terram Chananaei, Hetthaei et Amorraeiet Pherezaei et Iebusaei et Gergesaei,nempe ut dares semini eius;et implesti verba tua,quoniam iustus es.
NEH|9|9|Et vidisti afflictionem patrum nostrorum in Aegyptoclamoremque eorum audisti iuxta mare Rubrum.
NEH|9|10|Et dedisti signa atque portenta in pharaoneet in universis servis eius et in omni populo terrae illius;cognovisti enim quia superbe egerant contra eos,et fecisti tibi nomen, sicut et in hac die.
NEH|9|11|Et mare divisisti ante eos,et transierunt per medium maris in sicco;persecutores autem eorum proiecisti in profundum,quasi lapidem in aquas validas.
NEH|9|12|Et in columna nubis ductor eorum fuisti per diemet in columna ignis per noctem,ut illuminaret eis viam, per quam ingrediebantur.
NEH|9|13|Ad montem quoque Sinai descendistiet locutus es cum eis de caelo;et dedisti eis iudicia rectaet legem rectam, mandata et praecepta bona.
NEH|9|14|Et sabbatum sanctificatum tuum ostendisti eiset praecepta et mandata et legem praecepisti eisin manu Moysi servi tui.
NEH|9|15|Panem quoque de caelo dedisti eis in fame eorumet aquam de petra eduxisti eis in siti eorum;et dixisti eis, ut ingrederentur et possiderent terram,super quam levasti manum tuam, ut traderes eis.
NEH|9|16|Ipsi vero patres nostri superbe egeruntet induraverunt cervices suas et non audierunt mandata tua.
NEH|9|17|Et noluerunt audireet non sunt recordati mirabilium tuorum, quae feceras eis,et induraverunt cervices suaset posuerunt caput suum,ut reverterentur ad servitutem suam in Aegyptum.Tu autem Deus propitius, clemens et misericors,longanimis et multae miserationis, non dereliquisti eos.
NEH|9|18|Et quidem, cum fecissent sibi vitulum conflatilemet dixissent: "Iste est Deus tuus,qui eduxit te de Aegypto"feceruntque blasphemias magnas;
NEH|9|19|tu autem in misericordiis tuis multisnon dimisisti eos in deserto:columna nubis non recessit ab eis per diem,ut duceret eos in viam;et columna ignis per noctem,ut illuminaret eis iter, per quod ingrederentur.
NEH|9|20|Et spiritum tuum bonum dedisti, qui doceret eos,et manna tuum non prohibuisti ab ore eorumet aquam dedisti eis in siti eorum.
NEH|9|21|Quadraginta annis pavisti eos in deserto,nihilque eis defuit;vestimenta eorum non inveteraverunt,et pedes eorum non intumuerunt.
NEH|9|22|Et dedisti eis regna et populoset partitus es eis sortes;et possederunt terram Sehon et terram regis Hesebonet terram Og regis Basan.
NEH|9|23|Et multiplicasti filios eorum sicut stellas caeli;et adduxisti eos ad terram, de qua dixeras patribus eorum,ut ingrederentur et possiderent.
NEH|9|24|Et venerunt filii et possederunt terram,et humiliasti coram eis habitatores terrae Chananaeos;et dedisti eos in manu eorumet reges eorum et populos terrae,ut facerent eis, sicut placebat illis.
NEH|9|25|Ceperunt itaque urbes munitas et humum pinguem;et possederunt domos plenas cunctis bonis,cisternas ab aliis fabricatas, vineas et olivetaet ligna pomifera multa.Et comederunt et saturati sunt et impinguati suntet delectati sunt in bonitate tua magna.
NEH|9|26|Vexaverunt autem te et rebellaverunt contra teet proiecerunt legem tuam post terga sua;et prophetas tuos occiderunt,qui contestabantur eos, ut reverterentur ad te;feceruntque blasphemias grandes.
NEH|9|27|Et dedisti eos in manu hostium suorum,et afflixerunt eos;et in tempore tribulationis suae clamaverunt ad te,et tu de caelo audistiet secundum miserationes tuas multas dedisti eis salvatores,qui salvarent eos da manu hostium suorum.
NEH|9|28|Cumque requievissent, reversi sunt,ut facerent malum in conspectu tuo;et dereliquisti eos in manu inimicorum suorum,et dominati sunt eis.Conversique sunt et clamaverunt ad te;tu autem de caelo exaudistiet liberasti eos in misericordiis tuis multis vicibus.
NEH|9|29|Et contestatus es eos, ut reduceres eos ad legem tuam;ipsi vero superbe egerunt et non audierunt mandata tuaet in iudicia tua peccaverunt, quae si fecerit homo, vivet in eis, et dederunt umerum rebellemet cervicem suam induraverunt nec audierunt.
NEH|9|30|Et pepercisti eis annos multoset contestatus es eos in spiritu tuoper manum prophetarum tuorum, et non audierunt;et tradidisti eos in manu populorum terrarum.
NEH|9|31|In misericordiis autem tuis plurimisnon fecisti eos in consumptionemnec dereliquisti eos;quoniam Deus misericors et clemens es tu.
NEH|9|32|Nunc itaque, Deus noster magne, fortis et terribilis,custodiens pactum et misericordiam,ne parvipendas omnem laborem,qui invenit nos, reges nostros et principes nostroset sacerdotes nostros et prophetas nostroset patres nostros et omnem populum tuuma diebus regum Assyriae usque in diem hanc.
NEH|9|33|Et tu iustus es in omnibus, quae venerunt super nos,quia recte fecisti,nos autem impie egimus.
NEH|9|34|Reges nostri, principes nostri, sacerdotes nostri et patres nostrinon fecerunt legem tuamet non attenderunt mandata tua et testimonia tua,quae testificatus es in eis.
NEH|9|35|Et ipsi in regnis suis et in bonitate tua multa, quam dederas eis,et in terra latissima et pingui,quam tradideras in conspectu eorum,non servierunt tibi nec reversi sunt a studiis suis pessimis.
NEH|9|36|Ecce nos ipsi hodie servi sumus;et in terra, quam dedisti patribus nostris,ut comederent fructum eius et bona eius, nos ipsi servi sumus.
NEH|9|37|Et fruges eius multiplicantur regibus,quos posuisti super nos propter peccata nostra,et corporibus nostris dominantur et iumentis nostrissecundum voluntatem suam,et in tribulatione magna sumus ".
NEH|10|1|" Super omnibus ergo his nos ipsi percutimus foedus et scribimus, et signant principes nostri, Levitae nostri et sacerdotes nostri ".
NEH|10|2|Signatores autem fuerunt: Nehemias praepositus, filius Hachaliae, et Sedecias,
NEH|10|3|Saraias, Azarias, Ieremias,
NEH|10|4|Phassur, Amarias, Melchias,
NEH|10|5|Hattus, Sebania, Melluch,
NEH|10|6|Harim, Meremoth, Abdias,
NEH|10|7|Daniel, Genthon, Baruch,
NEH|10|8|Mosollam, Abia, Miamin,
NEH|10|9|Maazia, Belgai, Semeia; hi sacerdotes.
NEH|10|10|Porro Levitae: Iesua filius Azaniae, Bennui de filiis Henadad, Cadmihel
NEH|10|11|et fratres eorum Sebania, Hodia, Celita, Phalaia, Hanan,
NEH|10|12|Micha, Rohob, Hasabia,
NEH|10|13|Zacchur, Serebia, Sebania,
NEH|10|14|Hodia, Bani, Baninu.
NEH|10|15|Capita populi: Pharos, Phahathmoab, Elam, Zethua, Bani,
NEH|10|16|Bunni, Azgad, Bebai,
NEH|10|17|Adonia, Beguai, Adin,
NEH|10|18|Ater, Ezechia, Azur,
NEH|10|19|Hodia, Hasum, Besai,
NEH|10|20|Hareph, Anathoth, Nebai,
NEH|10|21|Megphias, Mosollam, Hezir,
NEH|10|22|Mesezabel, Sadoc, Ieddua,
NEH|10|23|Pheltia, Hanan, Anaia,
NEH|10|24|Osee, Hanania, Hassub,
NEH|10|25|Alohes, Phalea, Sobec,
NEH|10|26|Rehum, Hasabna, Maasia,
NEH|10|27|Ahia, Hanan, Anan,
NEH|10|28|Melluch, Harim, Baana.
NEH|10|29|Et reliqui de populo, sacerdotes, Levitae, ianitores et cantores, oblati et omnes, qui se separaverunt de populis terrarum ad legem Dei, uxores eorum, filii eorum et filiae eorum, omnes, qui poterant sapere,
NEH|10|30|adhaeserunt fratribus suis optimatibus pollicentes et iurantes, ut ambularent in lege Dei, quam dederat in manu Moysi servi Dei, et ut facerent et custodirent universa mandata Domini Dei nostri et iudicia eius et praecepta eius,
NEH|10|31|et ut non daremus filias nostras populo terrae et filias eorum non acciperemus filiis nostris.
NEH|10|32|Et si populi terrae importaverint venalia et omnia cibaria per diem sabbati, ut vendant, non accipiemus ab eis in sabbato et in die sanctificato; et dimittemus annum septimum et omnem exactionem.
NEH|10|33|Et statuimus super nos praecepta, ut demus tertiam partem sicli per annum ad opus domus Dei nostri,
NEH|10|34|ad panes propositionis et ad oblationem sempiternam et in holocaustum sempiternum in sabbatis, in calendis, in sollemnitatibus et in sanctificata et in sacrificium pro peccato, ut expietur pro Israel, et in omnem usum domus Dei nostri.
NEH|10|35|Sortes ergo misimus super oblationem lignorum inter sacerdotes et Levitas et populum, ut inferrentur in domum Dei nostri per domos patrum nostrorum, in temporibus constitutis ab anno in annum, ut arderent super altare domini Dei nostri, sicut scriptum est in lege;
NEH|10|36|et ut afferremus primogenita terrae nostrae et primitiva universi fructus omnis ligni ab anno in annum in domo Domini,
NEH|10|37|et primitiva filiorum nostrorum et pecorum nostrorum, sicut scriptum est in lege, et primitiva boum nostrorum et ovium nostrarum, ut afferrentur in domum Dei nostri sacerdotibus, qui ministrant in domo Dei nostri;
NEH|10|38|et primitias ciborum nostrorum et libaminum nostrorum et poma omnis ligni, vindemiae quoque et olei, afferemus sacerdotibus ad gazophylacium Dei nostri, et decimam partem terrae nostrae Levitis. Ipsi Levitae decimas accipient ex omnibus civitatibus agriculturae nostrae.
NEH|10|39|Erit autem sacerdos filius Aaron cum Levitis in decimis Levitarum colligendis, et Levitae offerent decimam partem decimae in domo Dei nostri ad gazophylacium thesauri.
NEH|10|40|Ad gazophylacium enim deportabunt filii Israel et filii Levi primitias frumenti, vini et olei; et ibi erunt vasa sanctificata et sacerdotes, qui ministrabant, et ianitores et cantores. Et non dimittemus domum Dei nostri.
NEH|11|1|Habitaverunt autem princi pes populi in Ierusalem; reli qua vero plebs misit sortem, ut adducerent unum virum de decem ad habitandum in Ierusalem civitate sancta, novem vero partes in civitatibus.
NEH|11|2|Benedixit autem populus omnibus viris, qui se sponte obtulerant, ut habitarent in Ierusalem.
NEH|11|3|Hi sunt itaque principes provinciae, qui habitaverunt in Ierusalem et in civitatibus Iudae. Habitavit autem unusquisque in possessione sua, in urbibus suis, Israel, sacerdotes, Levitae, oblati et filii servorum Salomonis.
NEH|11|4|Et in Ierusalem habitaverunt de filiis Iudae et de filiis Beniamin. De filiis Iudae: Athaias filius Oziam filii Zachariae filii Amariae filii Saphatiae filii Malaleel, de filiis Phares;
NEH|11|5|et Maasia filius Baruch filius Cholhoza filius Hazia filius Adaia filius Ioiarib filius Zachariae filius Silonitis.
NEH|11|6|Omnes filii Phares, qui habitaverunt in Ierusalem, quadringenti sexaginta octo viri fortes.
NEH|11|7|Hi sunt autem filii Beniamin: Sallu filius Mosollam filius Ioed filius Phadaia filius Colaia filius Maasia filius Etheel filius Iesaia;
NEH|11|8|et fratres eius viri fortes, nongenti viginti octo.
NEH|11|9|Et Ioel filius Zechri praepositus eorum, et Iudas filius Asana super civitatem secundus.
NEH|11|10|Et de sacerdotibus: Iedaia filius Ioiarib filius
NEH|11|11|Saraia filius Helciae filius Mosollam filius Sadoc filius Meraioth filius Achitob princeps domus Dei;
NEH|11|12|et fratres eorum facientes opera templi, octingenti viginti duo. Et Adaia filius Ieroham filius Phelelia filius Amsi filius Zachariae filius Phassur filius Melchiae;
NEH|11|13|et fratres eius principes familiarum ducenti quadraginta duo. Et Amassai filius Azareel filius Ahazi filius Mosollamoth filius Emmer;
NEH|11|14|et fratres eorum potentes nimis, centum viginti octo; et praepositus eorum Zabdiel vir nobilis.
NEH|11|15|Et de Levitis: Semeia filius Hassub filius Ezricam filius Hasabia filius Bunni;
NEH|11|16|et Sabethai et Iozabad super omnia opera, quae erant forinsecus in domo Dei, de principibus Levitarum;
NEH|11|17|et Matthania filius Micha filius Zebedaei filius Asaph magister chori incohabat orationem; et Becbecia secundus de fratribus eius, et Abda filius Sammua filius Galal filius Idithun.
NEH|11|18|Omnes Levitae in civitate sancta ducenti octoginta quattuor.
NEH|11|19|Et ianitores: Accub, Telmon et fratres eorum, qui custodiebant ostia, centum septuaginta duo.
NEH|11|20|Et reliqui ex Israel sacerdotes et Levitae in universis civitatibus Iudae, unusquisque in possessione sua.
NEH|11|21|Et oblati habitabant in Ophel; et Siha et Gaspha super oblatos.
NEH|11|22|Et praefectus Levitarum in Ierusalem Ozi filius Bani filius Hasabiae filius Matthaniae filius Michae de filiis Asaph, cantores in ministerio domus Dei.
NEH|11|23|Praeceptum quippe regis super eos erat, et ordo in cantoribus per dies singulos.
NEH|11|24|Et Phethahia filius Mesezabel de filiis Zara filii Iudae, legatus regis in omni negotio populi.
NEH|11|25|Et in viculis per omnes regiones eorum, de filiis Iudae habitaverunt in Cariatharbe et in pagis eius et in Dibon et in pagis eius et in Cabseel et in viculis eius
NEH|11|26|et in Iesua et in Molada et in Bethpheleth
NEH|11|27|et in Asarsual et in Bersabee et in pagis eius
NEH|11|28|et in Siceleg et in Mochona et in pagis eius
NEH|11|29|et in Remmon et in Saraa et in Ierimoth,
NEH|11|30|Zanoa, Odollam et in villis earum, Lachis et regionibus eius et Azeca et pagis eius. Et habitaverunt a Bersabee usque ad vallem Ennom.
NEH|11|31|Filii autem Beniamin in Gabaa, Machmas et Hai et Bethel et pagis eius,
NEH|11|32|Anathoth, Nob, Anania,
NEH|11|33|Asor, Rama, Getthaim,
NEH|11|34|Hadid, Seboim et Neballat,
NEH|11|35|Lod et Ono et valle Artificum.
NEH|11|36|Et de Levitis portiones in Iuda et Beniamin.
NEH|12|1|Hi sunt autem sacerdotes et Levitae, qui ascenderunt cum Zorobabel filio Salathiel et Iesua: Saraia, Ieremias, Esdras,
NEH|12|2|Amaria, Melluch, Hattus,
NEH|12|3|Sechenias, Rehum, Meremoth,
NEH|12|4|Addo, Genthon, Abia,
NEH|12|5|Miamin, Maadia, Belga,
NEH|12|6|Semeia et Ioiarib, Iedaia,
NEH|12|7|Sallu, Amoc, Helcias, Iedaia. Isti principes sacerdotum et fratrum eorum in diebus Iesua.
NEH|12|8|Porro Levitae: Iesua, Bennui, Cadmihel, Serebia, Iuda, Matthanias, super hymnos ipse et fratres eius;
NEH|12|9|et Becbecia atque Hanni fratres eorum coram eis per vices suas.
NEH|12|10|Iesua autem genuit Ioachim, et Ioachim genuit Eliasib, et Eliasib genuit Ioiada,
NEH|12|11|et Ioiada genuit Ionathan, et Ionathan genuit Ieddua.
NEH|12|12|In diebus autem Ioachim erant sacerdotes principes familiarum: Saraiae Maraia, Ieremiae Hanania,
NEH|12|13|Esdrae Mosollam, Amariae Iohanan,
NEH|12|14|Milicho Ionathan, Sebaniae Ioseph,
NEH|12|15|Harim Edna, Meraioth Helci,
NEH|12|16|Adaiae Zacharia, Genthon Mosollam,
NEH|12|17|Abiae Zechri, Miamin Maadiae Phelti,
NEH|12|18|Belgae Sammua, Semeiae Ionathan,
NEH|12|19|Ioiarib Matthanai, Iedaiae Ozi,
NEH|12|20|Sellai Celai, Amoc Heber,
NEH|12|21|Helciae Hasabia, Iedaiae Nathanael.
NEH|12|22|Levitae in diebus Eliasib et Ioiada et Iohanan et Ieddua scripti principes familiarum et sacerdotes usque ad regnurn Darii Persae.
NEH|12|23|Filii Levi principes familiarum scripti in libro Chronicorum usque ad dies Ionathan filii Eliasib.
NEH|12|24|Et principes Levitarum Hasabia, Serebia, Iesua, Bennui et Cadmihel et fratres eorum coram eis, ut laudarent et confiterentur iuxta praeceptum David viri Dei per vices suas;
NEH|12|25|Matthania et Becbecia, Abdia, Mosollam, Telmon, Accub ianitores ad custodiam horreorum iuxta portas.
NEH|12|26|Hi in diebus Ioachim filii Iesua filii Iosedec et in diebus Nehemiae ducis et Esdrae sacerdotis scribaeque.
NEH|12|27|In dedicatione autem muri Ierusalem requisierunt Levitas de omnibus locis suis, ut adducerent eos in Ierusalem et facerent dedicationem in laetitia, in actione gratiarum et cantico et cymbalis, psalteriis et citharis.
NEH|12|28|Congregati sunt autem cantores de campestribus circa Ierusalem et de villis Netophathitarum
NEH|12|29|et de Bethgalgala et de regionibus Gabaa et Azmaveth, quoniam villas aedificaverunt sibi cantores in circuitu Ierusalem.
NEH|12|30|Et mundati sunt sacerdotes et Levitae et mundaverunt populum et portas et murum.
NEH|12|31|Ascendere autem feci principes Iudae super murum et statui duos magnos choros laudantium, quorum unus ivit ad dexteram super murum ad portam Sterquilinii.
NEH|12|32|Et ivit post eos Osaias et media pars principum Iudae
NEH|12|33|et Azarias, Esdras et Mosollam,
NEH|12|34|Iudas et Beniamin et Semeia et Ieremias.
NEH|12|35|Et de sacerdotibus cum tubis et Zacharias filius Ionathan filius Semeiae filius Matthaniae filius Michaiae filius Zacchur filius Asaph;
NEH|12|36|et fratres eius Semeia et Azareel, Malalai, Galalai, Maai, Nathanael et Iudas et Hanani cum musicis David viri Dei; et Esdras scriba ante eos et in porta Fontis.
NEH|12|37|Processerunt per gradus civitatis David in ascensu muri super domum David et usque ad portam Aquarum ad orientem.
NEH|12|38|Et chorus secundus gratias referentium ibat ex adverso, et ego post eum, et media pars populi super murum et super turrim Furnorum et usque ad murum latissimum
NEH|12|39|et super portam Ephraim et super portam Antiquam et super portam Piscium et turrim Hananeel et turrim Meah et usque ad portam Gregis; et steterunt in porta Custodiae.
NEH|12|40|Steteruntque duo chori laudantium in domo Dei, et ego et dimidia pars magistratuum mecum.
NEH|12|41|Et sacerdotes Eliachim, Maasia, Miamin, Michaia, Elioenai, Zacharia, Hanania in tubis;
NEH|12|42|et Maasia et Semeia et Eleazar et Ozi et Iohanan et Melchia et Elam et Ezer. Et clare cecinerunt cantores et Izrahia praepositus.
NEH|12|43|Et obtulerunt in die illa sacrificia magna et laetati sunt; Deus enim laetificaverat eos laetitia magna; sed et uxores eorum et liberi gavisi sunt, et audita est laetitia Ierusalem procul.
NEH|12|44|Praeposuerunt quoque in die illa viros super gazophylacia ad thesaurum, ad libamina et ad primitias et ad decimas, ut colligerent in ea de agris civitatum partes legitimas pro sacerdotibus et Levitis; quia laetificatus est Iuda in sacerdotibus et Levitis, qui adstiterunt
NEH|12|45|et servierunt in ministerio Dei sui et in ministerio purificationis simul cum cantoribus et ianitoribus iuxta praeceptum David et Salomonis filii eius;
NEH|12|46|quia in diebus David et Asaph ab exordio erant catervae cantorum et carmina laudis et actionis gratiarum Deo.
NEH|12|47|Et omnis Israel in diebus Zorobabel et in diebus Nehemiae dabant partes cantoribus et ianitoribus per dies singulos partem suam et partes consecrabant Levitis, et Levitae consecrabant filiis Aaron.
NEH|13|1|In die autem illo lectum est in volumine Moysi, audiente populo, et inventum est scriptum in eo quod non debeant introire Ammonites et Moabites in ecclesiam Dei usque in aeternum,
NEH|13|2|eo quod non occurrerint filiis Israel cum pane et aqua et conduxerint adversum eos Balaam ad maledicendum eis, et convertit Deus noster maledictionem in benedictionem.
NEH|13|3|Factum est autem, cum audissent legem, separaverunt omnem promiscuum ab Israel.
NEH|13|4|Ante hoc autem erat Eliasib sacerdos, qui fuerat praepositus in gazophylacio domus Dei nostri et proximus Thobiae;
NEH|13|5|fecerat ei gazophylacium grande, ubi antea reponebant munera et tus et vasa et decimam frumenti, vini et olei, partes Levitarum et cantorum et ianitorum et tributa sacerdotum.
NEH|13|6|In omnibus autem his non fui in Ierusalem, quia anno tricesimo secundo Artaxerxis regis Babylonis veni ad regem et in fine dierum rogavi, ut abirem a rege,
NEH|13|7|et veni in Ierusalem. Et intellexi malum, quod fecerat Eliasib Thobiae: fecerat enim ei thesaurum in vestibulis domus Dei.
NEH|13|8|Et malum mihi visum est valde, et proieci vasa domus Thobiae foras de gazophylacio;
NEH|13|9|praecepique, et emundaverunt gazophylacia, et rettuli ibi vasa domus Dei, oblationem et tus.
NEH|13|10|Et cognovi quod partes Levitarum non fuissent datae, et fugisset unusquisque in campum suum de Levitis et cantoribus, qui ministrabant.
NEH|13|11|Et egi causam adversus magistratus et dixi: " Quare dereliquimus domum Dei? ". Et congregavi eos et feci stare in stationibus suis.
NEH|13|12|Et omnis Iuda apportabat decimam frumenti, vini et olei in horrea.
NEH|13|13|Et constitui super horrea Selemiam sacerdotem et Sadoc scribam et Phadaiam de Levitis et iuxta eos Hanan filium Zacchur, filium Matthaniae, quoniam fideles comprobati sunt; et ipsi curam habebant distribuendi partes fratribus suis.
NEH|13|14|Memento mei, Deus meus, pro hoc; et ne deleas opera mea bona, quae feci in domo Dei mei et in ministeriis eius!
NEH|13|15|In diebus illis vidi in Iuda calcantes torcularia in sabbato, portantes acervos et onerantes super asinos vinum et uvas et ficus et omne onus et inferentes in Ierusalem die sabbati; et contestatus sum, quando vendebant cibaria.
NEH|13|16|Et ibi Tyrii habitaverunt in ea inferentes pisces et omnia venalia et vendebant in sabbatis filiis Iudae in Ierusalem.
NEH|13|17|Et obiurgavi optimates Iudae et dixi eis: " Quae est haec res mala, quam vos facitis, et profanatis diem sabbati?
NEH|13|18|Numquid non haec fecerunt patres nostri, et adduxit Deus noster super nos omne malum hoc et super civitatem hanc? Et vos additis iracundiam super Israel profanando sabbatum! ".
NEH|13|19|Factum est autem, cum obscuratae essent portae Ierusalem ante diem sabbati, dixi, et clauserunt ianuas; et praecepi, ut non aperirent eas usque post sabbatum. Et de pueris meis constitui super portas, ut nullus inferret onus in die sabbati.
NEH|13|20|Et manserunt negotiatores et vendentes universa venalia foris Ierusalem semel et bis.
NEH|13|21|Et contestatus sum eos et dixi eis: " Quare manetis ex adverso muri? Si iterum hoc feceritis, manum mittam in vos ". Itaque ex tempore illo non venerunt in sabbato.
NEH|13|22|Dixi quoque Levitis, ut mundarentur et venirent ad custodiendas portas et sanctificandam diem sabbati.Et pro hoc ergo memento mei, Deus meus, et parce mihi secundum multitudinem miserationum tuarum!
NEH|13|23|Sed et in diebus illis vidi Iudaeos, qui duxerant uxores Azotidas, Ammonitidas et Moabitidas.
NEH|13|24|Et filii eorum ex media parte loquebantur Azotice et nesciebant loqui Iudaice vel loquebantur iuxta linguam unius vel alterius populi.
NEH|13|25|Et obiurgavi eos et maledixi et cecidi quosdam ex eis et decalvavi eos; et adiuravi in Deo, ut non darent filias suas filiis eorum et non acciperent de filiabus eorum filiis suis et sibimetipsis dicens:
NEH|13|26|" Numquid non in huiuscemodi re peccavit Salomon rex Israel? Et certe in gentibus multis non erat rex similis ei, et dilectus Deo suo erat, et posuit eum Deus regem super omnem Israel; et ipsum ergo duxerunt ad peccatum mulieres alienigenae.
NEH|13|27|Numquid et vobis obsequentes faciemus omne malum grande hoc, ut praevaricemur in Deo nostro et ducamus uxores peregrinas? ".
NEH|13|28|Unus autem de filiis Ioiada filii Eliasib sacerdotis magni gener erat Sanaballat Horonites, quem fugavi a me.
NEH|13|29|Recordare, Domine Deus meus, adversum eos, qui polluunt sacerdotium et pactum sacerdotale et leviticum!
NEH|13|30|Igitur mundavi eos ab omnibus alienigenis et constitui ordines pro sacerdotibus et Levitis, unumquemque in ministerio suo,
NEH|13|31|et pro oblatione lignorum in temporibus constitutis et pro primitiis. Memento mei, Deus meus, in bonum.
