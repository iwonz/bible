JAS|1|1|上帝和主耶穌基督的僕人 雅各 問候散居在各處的十二個支派的人。
JAS|1|2|我的弟兄們，你們遭受各種試煉時，都要認為是大喜樂，
JAS|1|3|因為知道你們的信心經過考驗，就生忍耐。
JAS|1|4|但要讓忍耐發揮完全的功用，使你們能又完全又完整，一無所缺。
JAS|1|5|你們中間若有缺少智慧的，該求那厚賜與眾人又不斥責人的上帝，上帝必賜給他。
JAS|1|6|只要憑著信心求，一點也不疑惑；因為那疑惑的人，就像海中的波浪被風吹動翻騰。
JAS|1|7|這樣的人不要想從主那裏得到甚麼。
JAS|1|8|三心二意的人，在他一切所行的路上都搖擺不定。
JAS|1|9|卑微的弟兄要因高升而誇耀，
JAS|1|10|富足的卻要因被降卑而誇耀，因為富足的人要消逝，如同草上的花一樣。
JAS|1|11|太陽出來，熱風颳起，草就枯乾，花也凋謝，它美麗的樣子就消失了；那富足的人在他一生的奔波中也要這樣衰殘。
JAS|1|12|忍受試煉的人有福了，因為他經過考驗以後必得生命的冠冕，這是主應許給愛他之人的。
JAS|1|13|人被誘惑，不可說：「我是被上帝誘惑」；因為上帝是不被惡誘惑的，他也不誘惑人。
JAS|1|14|但每一個人被誘惑是因自己的私慾牽引而被誘惑的。
JAS|1|15|私慾既懷了胎，就生出罪來；罪既長成，就生出死來。
JAS|1|16|我親愛的弟兄們，不要被欺騙了。
JAS|1|17|各樣美善的恩澤和各樣完美的賞賜都是從上頭來的，從眾光之父那裏降下來的；在他並沒有改變，也沒有轉動的影兒。
JAS|1|18|他按自己的旨意，用真理的道生了我們，使我們在他所造的萬物中成為初熟的果子。
JAS|1|19|我親愛的弟兄們，你們要明白：你們每一個人要快快地聽，慢慢地說，慢慢地動怒，
JAS|1|20|因為人的怒氣並不能實現上帝的義。
JAS|1|21|所以，你們要除去一切的污穢和累積的惡毒，要存溫柔的心領受所栽種的道，就是能救你們靈魂的道。
JAS|1|22|但是，你們要作行道的人，不要只作聽道的人，自己欺騙自己。
JAS|1|23|因為只聽道而不行道的，就像人對著鏡子觀看自己本來的面目，
JAS|1|24|注視後，就離開，立刻忘了自己的相貌如何。
JAS|1|25|惟有查看那完美、使人自由的律法，並且時常遵守的，他不是聽了就忘，而是切實行出來，這樣的人在所行的事上必然蒙福。
JAS|1|26|若有人自以為虔誠，卻不勒住自己的舌頭，反欺騙自己的心，這人的虔誠是徒然的。
JAS|1|27|在上帝—我們的父面前，清潔沒有玷污的虔誠就是看顧在患難中的孤兒寡婦，並且保守自己不沾染世俗。
JAS|2|1|我的弟兄們，你們信奉我們榮耀的主耶穌基督，就不可按著外貌待人。
JAS|2|2|若有一個人戴著金戒指，穿著華麗的衣服，進入你們的會堂，又有一個窮人穿著骯髒的衣服也進去，
JAS|2|3|而你們只看重那穿華麗衣服的人，說：「請坐在這裏」，又對那窮人說：「你站在那裏」，或「坐在我腳凳旁」；
JAS|2|4|這豈不是你們偏心待人，用惡意評斷人嗎？
JAS|2|5|我親愛的弟兄們，請聽，上帝豈不是揀選了世上的貧窮人，使他們在信心上富足，並承受他所應許給那些愛他之人的國嗎？
JAS|2|6|你們卻羞辱貧窮的人。欺壓你們，拉你們到公堂去的，不就是這些富有的人嗎？
JAS|2|7|毀謗為你們求告時所奉的尊名的，不就是他們嗎？
JAS|2|8|經上記著：「要愛鄰 如己」，你們若切實守這至尊的律法，你們就做得很好。
JAS|2|9|但你們若按外貌待人就是犯罪，是被律法定為犯法的。
JAS|2|10|因為凡遵守全部律法的，只違背了一條就是違犯了所有的律法。
JAS|2|11|原來那說「不可姦淫」的，也說「不可殺人」。你就是不姦淫，卻殺人，也是成為違犯律法的。
JAS|2|12|既然你們要按使人自由的律法受審判，就要照這律法說話行事。
JAS|2|13|因為對那不憐憫人的，他們要受沒有憐憫的審判；憐憫勝過審判。
JAS|2|14|我的弟兄們，若有人說自己有信心，卻沒有行為，有甚麼益處呢？這信心能救他嗎？
JAS|2|15|若是弟兄或是姊妹沒有衣服穿，又缺少日用的飲食；
JAS|2|16|你們中間有人對他們說：「平平安安地去吧！願你們穿得暖，吃得飽」，卻不給他們身體所需要的，這有甚麼益處呢？
JAS|2|17|信心也是這樣，若沒有行為是死的。
JAS|2|18|但是有人會說：「你有信心，我有行為。」把你沒有行為的信心給我看，我就藉著我的行為把我的信心給你看。
JAS|2|19|你信上帝只有一位，你信得很好；連鬼魔也信，且怕得發抖。
JAS|2|20|你這虛浮的人哪，你願意知道沒有行為的信心是沒有用的嗎？
JAS|2|21|我們的祖宗 亞伯拉罕 把他兒子 以撒 獻在壇上，豈不是因行為得稱義嗎？
JAS|2|22|可見信心是與他的行為相輔並行，而且信心是因著行為才得以成全的。
JAS|2|23|這正應驗了經上所說：「 亞伯拉罕 信了上帝，這就算他為義」；他又得稱為上帝的朋友。
JAS|2|24|這樣看來，人稱義是因著行為，不是單因著信。
JAS|2|25|同樣，妓女 喇合 接待使者，又放他們從另一條路出去，不也是因行為稱義嗎？
JAS|2|26|所以，就如身體沒有靈魂是死的，信心沒有行為也是死的。
JAS|3|1|我的弟兄們，不要許多人做教師，因為你們知道，我們做教師的要接受更嚴厲的審判。
JAS|3|2|原來我們在許多事上都有過失；若有人在言語上沒有過失，他就是完全的人，也能勒住自己的全身。
JAS|3|3|我們若把嚼環放在馬嘴裏使牠們馴服，就能控制牠們的全身。
JAS|3|4|再看船隻，雖然甚大，又被強風猛吹，只用小小的舵就隨著掌舵的意思轉動。
JAS|3|5|同樣，舌頭是小肢體，卻能說大話。 看哪，最小的火能點燃最大的樹林。
JAS|3|6|舌頭就是火。在我們百體中，舌頭是個不義的世界，能玷污全身，也能燒燬生命的輪子，而且是被地獄的火點燃的。
JAS|3|7|各類的走獸、飛禽、爬蟲、水族，本來都可以制伏，也已經被人制伏了；
JAS|3|8|惟獨舌頭沒有人能制伏，是永不靜止的邪惡，充滿了害死人的毒氣。
JAS|3|9|我們用舌頭頌讚我們的主—我們的天父，又用舌頭詛咒照著上帝形像被造的人。
JAS|3|10|頌讚和詛咒從同一個口出來。我的弟兄們，這是不應該的。
JAS|3|11|泉源能從一個出口發出甜苦兩樣的水嗎？
JAS|3|12|我的弟兄們，無花果樹能生橄欖嗎？葡萄樹能結無花果嗎？鹹水也不能流出甜水來。
JAS|3|13|你們中間誰是有智慧有見識的呢？他就當在智慧的溫柔上顯出他的善行來。
JAS|3|14|你們心裏若懷著惡毒的嫉妒和自私，就不可自誇，不可說謊話抵擋真理。
JAS|3|15|這樣的智慧不是從上頭下來的，而是屬地上的，屬情慾的，屬鬼魔的。
JAS|3|16|在何處有嫉妒、自私，在何處就有動亂和各樣的壞事。
JAS|3|17|惟獨從上頭來的智慧，先是清潔，後是和平、溫良、柔順，滿有憐憫和美善的果子，沒有偏私，沒有虛偽。
JAS|3|18|正義的果實是為促進和平的人用和平栽種出來的。
JAS|4|1|你們中間的衝突是哪裏來的？爭執是哪裏來的？不是從你們肢體中交戰著的私慾來的嗎？
JAS|4|2|你們貪戀，得不著就殺人；你們嫉妒，不能得手就起爭執和衝突；你們得不著，是因為你們不求。
JAS|4|3|你們求也得不著，是因為你們妄求，為了要浪費在你們的宴樂中。
JAS|4|4|你們這些淫亂的人哪，豈不知道與世俗為友就是與上帝為敵嗎？所以，凡想要與世俗為友的，就是與上帝為敵了。
JAS|4|5|經上說：「上帝愛安置在我們裏面的靈，愛到嫉妒的地步。」 你們以為這話是徒然的嗎？
JAS|4|6|但是他賜更多的恩典，正如經上說： 「上帝抵擋驕傲的人， 但賜恩給謙卑的人。」
JAS|4|7|所以，要順服上帝。要抵擋魔鬼，魔鬼就必逃避你們；
JAS|4|8|要親近上帝，上帝就必親近你們。有罪的人哪，要潔淨你們的手！心懷二意的人哪，要清潔你們的心！
JAS|4|9|你們要愁苦，悲哀，哭泣；要將歡笑變為悲哀，歡樂變為愁悶。
JAS|4|10|要在主面前謙卑，他就使你們高升。
JAS|4|11|弟兄們，不可彼此詆毀。詆毀弟兄或評斷弟兄的人，就是詆毀律法，評斷律法；你若評斷律法，就不是遵行律法，而是評斷者了。
JAS|4|12|立法者和審判者只有一位；他就是那能拯救人也能毀滅人的。你是誰，竟敢評斷你的鄰舍！
JAS|4|13|注意！有人說：「今天或明天我們要往某城去，在那裏住一年，做買賣賺錢。」
JAS|4|14|其實明天如何，你們還不知道。你們的生命是甚麼呢？你們 原來是一片雲霧，出現片刻就不見了。
JAS|4|15|你們倒應當說：「主若願意，我們就能活著，也可以做這事或那事。」
JAS|4|16|現今你們竟然狂傲自誇；凡這樣的自誇都是邪惡的。
JAS|4|17|所以，人若知道該行善而不去行，這就是他的罪了。
JAS|5|1|注意！你們這些富足人哪，要為將要臨到你們身上的災難哭泣、號咷。
JAS|5|2|你們的財物腐爛了，你們的衣服被蟲子蛀了。
JAS|5|3|你們的金銀都生銹了；這銹要證明你們的不是，又要像火一樣吞吃你們的肉。你們在這末世只知道積蓄錢財。
JAS|5|4|工人給你們收割莊稼，你們剋扣他們的工錢；這工錢在喊冤，而且收割工人的冤聲已經進入萬軍之主的耳朵了。
JAS|5|5|你們在地上享奢華宴樂，把自己養肥了，等候宰殺的日子。
JAS|5|6|你們定了義人的罪，把他殺害，他沒有抵抗你們。
JAS|5|7|所以弟兄們，你們要忍耐，直到主來。看哪，農夫等候著地裏寶貴的出產，耐心地等到它得了秋霖春雨。
JAS|5|8|你們也要忍耐，堅固你們的心，因為主來的日子近了。
JAS|5|9|弟兄們，你們不要彼此埋怨，免得受審判。看哪，審判的主站在門口了。
JAS|5|10|弟兄們，你們要把那先前奉主名說話的眾先知作能受苦、能忍耐的榜樣。
JAS|5|11|看哪，那些忍耐的人，我們稱他們是有福的。你們聽見過 約伯 的忍耐，也看見主給他的結局，知道主是充滿憐憫和慈悲的。
JAS|5|12|我的弟兄們，最要緊的是不可起誓；不可指著天起誓，也不可指著地起誓，任何誓都不可起。你們說話，是，就說是；不是，就說不是，免得你們落在審判之下。
JAS|5|13|你們中間若有人受苦，他該禱告；有人喜樂，他該歌頌。
JAS|5|14|你們中間若有人病了，他該請教會的長老們來為他禱告，奉主的名為他抹油。
JAS|5|15|出於信心的祈禱必能救那病人，主必叫他起來；他若犯了罪，也必蒙赦免。
JAS|5|16|所以，你們要彼此認罪，互相代求，使你們得醫治。義人祈禱所發的力量是大有功效的。
JAS|5|17|以利亞 與我們是同樣性情的人，他懇切地祈求不要下雨，地上就三年六個月沒有下雨。
JAS|5|18|他又禱告，天就降下雨來，地就有了出產。
JAS|5|19|我的弟兄們，你們中間若有人迷失了真理而有人使他回轉，
JAS|5|20|這人該知道，使一個罪人從迷途中回轉，會從死亡中把他的靈魂救回來，而且遮蓋許多的罪。
