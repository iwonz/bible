1PET|1|1|Peter, an apostle of Jesus Christ, to the strangers scattered throughout Pontus, Galatia, Cappadocia, Asia, and Bithynia,
1PET|1|2|Elect according to the foreknowledge of God the Father, through sanctification of the Spirit, unto obedience and sprinkling of the blood of Jesus Christ: Grace unto you, and peace, be multiplied.
1PET|1|3|Blessed be the God and Father of our Lord Jesus Christ, which according to his abundant mercy hath begotten us again unto a lively hope by the resurrection of Jesus Christ from the dead,
1PET|1|4|To an inheritance incorruptible, and undefiled, and that fadeth not away, reserved in heaven for you,
1PET|1|5|Who are kept by the power of God through faith unto salvation ready to be revealed in the last time.
1PET|1|6|Wherein ye greatly rejoice, though now for a season, if need be, ye are in heaviness through manifold temptations:
1PET|1|7|That the trial of your faith, being much more precious than of gold that perisheth, though it be tried with fire, might be found unto praise and honour and glory at the appearing of Jesus Christ:
1PET|1|8|Whom having not seen, ye love; in whom, though now ye see him not, yet believing, ye rejoice with joy unspeakable and full of glory:
1PET|1|9|Receiving the end of your faith, even the salvation of your souls.
1PET|1|10|Of which salvation the prophets have enquired and searched diligently, who prophesied of the grace that should come unto you:
1PET|1|11|Searching what, or what manner of time the Spirit of Christ which was in them did signify, when it testified beforehand the sufferings of Christ, and the glory that should follow.
1PET|1|12|Unto whom it was revealed, that not unto themselves, but unto us they did minister the things, which are now reported unto you by them that have preached the gospel unto you with the Holy Ghost sent down from heaven; which things the angels desire to look into.
1PET|1|13|Wherefore gird up the loins of your mind, be sober, and hope to the end for the grace that is to be brought unto you at the revelation of Jesus Christ;
1PET|1|14|As obedient children, not fashioning yourselves according to the former lusts in your ignorance:
1PET|1|15|But as he which hath called you is holy, so be ye holy in all manner of conversation;
1PET|1|16|Because it is written, Be ye holy; for I am holy.
1PET|1|17|And if ye call on the Father, who without respect of persons judgeth according to every man's work, pass the time of your sojourning here in fear:
1PET|1|18|Forasmuch as ye know that ye were not redeemed with corruptible things, as silver and gold, from your vain conversation received by tradition from your fathers;
1PET|1|19|But with the precious blood of Christ, as of a lamb without blemish and without spot:
1PET|1|20|Who verily was foreordained before the foundation of the world, but was manifest in these last times for you,
1PET|1|21|Who by him do believe in God, that raised him up from the dead, and gave him glory; that your faith and hope might be in God.
1PET|1|22|Seeing ye have purified your souls in obeying the truth through the Spirit unto unfeigned love of the brethren, see that ye love one another with a pure heart fervently:
1PET|1|23|Being born again, not of corruptible seed, but of incorruptible, by the word of God, which liveth and abideth for ever.
1PET|1|24|For all flesh is as grass, and all the glory of man as the flower of grass. The grass withereth, and the flower thereof falleth away:
1PET|1|25|But the word of the Lord endureth for ever. And this is the word which by the gospel is preached unto you.
1PET|2|1|Wherefore laying aside all malice, and all guile, and hypocrisies, and envies, all evil speakings,
1PET|2|2|As newborn babes, desire the sincere milk of the word, that ye may grow thereby:
1PET|2|3|If so be ye have tasted that the Lord is gracious.
1PET|2|4|To whom coming, as unto a living stone, disallowed indeed of men, but chosen of God, and precious,
1PET|2|5|Ye also, as lively stones, are built up a spiritual house, an holy priesthood, to offer up spiritual sacrifices, acceptable to God by Jesus Christ.
1PET|2|6|Wherefore also it is contained in the scripture, Behold, I lay in Sion a chief corner stone, elect, precious: and he that believeth on him shall not be confounded.
1PET|2|7|Unto you therefore which believe he is precious: but unto them which be disobedient, the stone which the builders disallowed, the same is made the head of the corner,
1PET|2|8|And a stone of stumbling, and a rock of offence, even to them which stumble at the word, being disobedient: whereunto also they were appointed.
1PET|2|9|But ye are a chosen generation, a royal priesthood, an holy nation, a peculiar people; that ye should shew forth the praises of him who hath called you out of darkness into his marvellous light;
1PET|2|10|Which in time past were not a people, but are now the people of God: which had not obtained mercy, but now have obtained mercy.
1PET|2|11|Dearly beloved, I beseech you as strangers and pilgrims, abstain from fleshly lusts, which war against the soul;
1PET|2|12|Having your conversation honest among the Gentiles: that, whereas they speak against you as evildoers, they may by your good works, which they shall behold, glorify God in the day of visitation.
1PET|2|13|Submit yourselves to every ordinance of man for the Lord's sake: whether it be to the king, as supreme;
1PET|2|14|Or unto governors, as unto them that are sent by him for the punishment of evildoers, and for the praise of them that do well.
1PET|2|15|For so is the will of God, that with well doing ye may put to silence the ignorance of foolish men:
1PET|2|16|As free, and not using your liberty for a cloke of maliciousness, but as the servants of God.
1PET|2|17|Honour all men. Love the brotherhood. Fear God. Honour the king.
1PET|2|18|Servants, be subject to your masters with all fear; not only to the good and gentle, but also to the froward.
1PET|2|19|For this is thankworthy, if a man for conscience toward God endure grief, suffering wrongfully.
1PET|2|20|For what glory is it, if, when ye be buffeted for your faults, ye shall take it patiently? but if, when ye do well, and suffer for it, ye take it patiently, this is acceptable with God.
1PET|2|21|For even hereunto were ye called: because Christ also suffered for us, leaving us an example, that ye should follow his steps:
1PET|2|22|Who did no sin, neither was guile found in his mouth:
1PET|2|23|Who, when he was reviled, reviled not again; when he suffered, he threatened not; but committed himself to him that judgeth righteously:
1PET|2|24|Who his own self bare our sins in his own body on the tree, that we, being dead to sins, should live unto righteousness: by whose stripes ye were healed.
1PET|2|25|For ye were as sheep going astray; but are now returned unto the Shepherd and Bishop of your souls.
1PET|3|1|Likewise, ye wives, be in subjection to your own husbands; that, if any obey not the word, they also may without the word be won by the conversation of the wives;
1PET|3|2|While they behold your chaste conversation coupled with fear.
1PET|3|3|Whose adorning let it not be that outward adorning of plaiting the hair, and of wearing of gold, or of putting on of apparel;
1PET|3|4|But let it be the hidden man of the heart, in that which is not corruptible, even the ornament of a meek and quiet spirit, which is in the sight of God of great price.
1PET|3|5|For after this manner in the old time the holy women also, who trusted in God, adorned themselves, being in subjection unto their own husbands:
1PET|3|6|Even as Sara obeyed Abraham, calling him lord: whose daughters ye are, as long as ye do well, and are not afraid with any amazement.
1PET|3|7|Likewise, ye husbands, dwell with them according to knowledge, giving honour unto the wife, as unto the weaker vessel, and as being heirs together of the grace of life; that your prayers be not hindered.
1PET|3|8|Finally, be ye all of one mind, having compassion one of another, love as brethren, be pitiful, be courteous:
1PET|3|9|Not rendering evil for evil, or railing for railing: but contrariwise blessing; knowing that ye are thereunto called, that ye should inherit a blessing.
1PET|3|10|For he that will love life, and see good days, let him refrain his tongue from evil, and his lips that they speak no guile:
1PET|3|11|Let him eschew evil, and do good; let him seek peace, and ensue it.
1PET|3|12|For the eyes of the Lord are over the righteous, and his ears are open unto their prayers: but the face of the Lord is against them that do evil.
1PET|3|13|And who is he that will harm you, if ye be followers of that which is good?
1PET|3|14|But and if ye suffer for righteousness' sake, happy are ye: and be not afraid of their terror, neither be troubled;
1PET|3|15|But sanctify the Lord God in your hearts: and be ready always to give an answer to every man that asketh you a reason of the hope that is in you with meekness and fear:
1PET|3|16|Having a good conscience; that, whereas they speak evil of you, as of evildoers, they may be ashamed that falsely accuse your good conversation in Christ.
1PET|3|17|For it is better, if the will of God be so, that ye suffer for well doing, than for evil doing.
1PET|3|18|For Christ also hath once suffered for sins, the just for the unjust, that he might bring us to God, being put to death in the flesh, but quickened by the Spirit:
1PET|3|19|By which also he went and preached unto the spirits in prison;
1PET|3|20|Which sometime were disobedient, when once the longsuffering of God waited in the days of Noah, while the ark was a preparing, wherein few, that is, eight souls were saved by water.
1PET|3|21|The like figure whereunto even baptism doth also now save us (not the putting away of the filth of the flesh, but the answer of a good conscience toward God,) by the resurrection of Jesus Christ:
1PET|3|22|Who is gone into heaven, and is on the right hand of God; angels and authorities and powers being made subject unto him.
1PET|4|1|Forasmuch then as Christ hath suffered for us in the flesh, arm yourselves likewise with the same mind: for he that hath suffered in the flesh hath ceased from sin;
1PET|4|2|That he no longer should live the rest of his time in the flesh to the lusts of men, but to the will of God.
1PET|4|3|For the time past of our life may suffice us to have wrought the will of the Gentiles, when we walked in lasciviousness, lusts, excess of wine, revellings, banquetings, and abominable idolatries:
1PET|4|4|Wherein they think it strange that ye run not with them to the same excess of riot, speaking evil of you:
1PET|4|5|Who shall give account to him that is ready to judge the quick and the dead.
1PET|4|6|For for this cause was the gospel preached also to them that are dead, that they might be judged according to men in the flesh, but live according to God in the spirit.
1PET|4|7|But the end of all things is at hand: be ye therefore sober, and watch unto prayer.
1PET|4|8|And above all things have fervent charity among yourselves: for charity shall cover the multitude of sins.
1PET|4|9|Use hospitality one to another without grudging.
1PET|4|10|As every man hath received the gift, even so minister the same one to another, as good stewards of the manifold grace of God.
1PET|4|11|If any man speak, let him speak as the oracles of God; if any man minister, let him do it as of the ability which God giveth: that God in all things may be glorified through Jesus Christ, to whom be praise and dominion for ever and ever. Amen.
1PET|4|12|Beloved, think it not strange concerning the fiery trial which is to try you, as though some strange thing happened unto you:
1PET|4|13|But rejoice, inasmuch as ye are partakers of Christ's sufferings; that, when his glory shall be revealed, ye may be glad also with exceeding joy.
1PET|4|14|If ye be reproached for the name of Christ, happy are ye; for the spirit of glory and of God resteth upon you: on their part he is evil spoken of, but on your part he is glorified.
1PET|4|15|But let none of you suffer as a murderer, or as a thief, or as an evildoer, or as a busybody in other men's matters.
1PET|4|16|Yet if any man suffer as a Christian, let him not be ashamed; but let him glorify God on this behalf.
1PET|4|17|For the time is come that judgment must begin at the house of God: and if it first begin at us, what shall the end be of them that obey not the gospel of God?
1PET|4|18|And if the righteous scarcely be saved, where shall the ungodly and the sinner appear?
1PET|4|19|Wherefore let them that suffer according to the will of God commit the keeping of their souls to him in well doing, as unto a faithful Creator.
1PET|5|1|The elders which are among you I exhort, who am also an elder, and a witness of the sufferings of Christ, and also a partaker of the glory that shall be revealed:
1PET|5|2|Feed the flock of God which is among you, taking the oversight thereof, not by constraint, but willingly; not for filthy lucre, but of a ready mind;
1PET|5|3|Neither as being lords over God's heritage, but being ensamples to the flock.
1PET|5|4|And when the chief Shepherd shall appear, ye shall receive a crown of glory that fadeth not away.
1PET|5|5|Likewise, ye younger, submit yourselves unto the elder. Yea, all of you be subject one to another, and be clothed with humility: for God resisteth the proud, and giveth grace to the humble.
1PET|5|6|Humble yourselves therefore under the mighty hand of God, that he may exalt you in due time:
1PET|5|7|Casting all your care upon him; for he careth for you.
1PET|5|8|Be sober, be vigilant; because your adversary the devil, as a roaring lion, walketh about, seeking whom he may devour:
1PET|5|9|Whom resist stedfast in the faith, knowing that the same afflictions are accomplished in your brethren that are in the world.
1PET|5|10|But the God of all grace, who hath called us unto his eternal glory by Christ Jesus, after that ye have suffered a while, make you perfect, stablish, strengthen, settle you.
1PET|5|11|To him be glory and dominion for ever and ever. Amen.
1PET|5|12|By Silvanus, a faithful brother unto you, as I suppose, I have written briefly, exhorting, and testifying that this is the true grace of God wherein ye stand.
1PET|5|13|The church that is at Babylon, elected together with you, saluteth you; and so doth Marcus my son.
1PET|5|14|Greet ye one another with a kiss of charity. Peace be with you all that are in Christ Jesus. Amen.
