PHLM|1|1|为基督耶稣被囚的 保罗 ，同弟兄 提摩太 ，写信给我们所亲爱的同工 腓利门 、
PHLM|1|2|亚腓亚 姊妹，和我们的战友 亚基布 ，以及在你家里的教会。
PHLM|1|3|愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
PHLM|1|4|我在祷告中记念你的时候，常为你感谢我的上帝，
PHLM|1|5|因听说你对众圣徒的爱心，和你对主耶稣的信心。
PHLM|1|6|愿你与人分享信心的时候，能产生功效，让人知道我们 所行的各样善事都是为基督做的。
PHLM|1|7|弟兄啊，由于你的爱心，我得到极大的快乐和安慰，因为众圣徒的心从你得到舒畅。
PHLM|1|8|虽然我靠着基督能放胆吩咐你做该做的事，
PHLM|1|9|可是像我这上了年纪的 保罗 ，现在又是为基督耶稣被囚的，宁可凭着爱心求你，
PHLM|1|10|就是为我在捆锁中所生的儿子 阿尼西谋 求你。
PHLM|1|11|从前他与你没有益处，但如今与你我都有益处。
PHLM|1|12|我现在打发他回到你那里去，他是我心肝。
PHLM|1|13|我本来有意将他留下，在我为福音所受的捆锁中替你伺候我。
PHLM|1|14|但不知道你的意见，我不愿意这样做，好使你的善行不是出于勉强，而是出于自愿。
PHLM|1|15|他暂时离开你，也许是要让你永远得着他，
PHLM|1|16|不再是奴隶，而是高过奴隶，是亲爱的弟兄；对我确实如此，何况对你呢！无论在肉身或在主里更是如此。
PHLM|1|17|所以，你若以我为同伴，就接纳他，如同接纳我一样。
PHLM|1|18|他若亏负你，或欠你什么，都算在我的账上吧，
PHLM|1|19|我必偿还。这是我— 保罗 亲笔写的。我并不用对你说，甚至你自己也亏欠我呢！
PHLM|1|20|弟兄啊，希望你使我在主里因你得益处，让我的心在基督里得到舒畅。
PHLM|1|21|我写信给你，深信你必顺服，知道你所要做的，必过于我所说的。
PHLM|1|22|此外，还请给我预备住处，因为我盼望藉着你们的祷告，必蒙恩回到你们那里去。
PHLM|1|23|为基督耶稣与我一同坐监的 以巴弗 问候你。
PHLM|1|24|我的同工 马可 、 亚里达古 、 底马 、 路加 也都问候你。
PHLM|1|25|愿 主耶稣基督的恩与你们的灵同在。
