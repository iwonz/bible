JOB|1|1|Был человек в земле Уц, имя его Иов; и был человек этот непорочен, справедлив и богобоязнен и удалялся от зла.
JOB|1|2|И родились у него семь сыновей и три дочери.
JOB|1|3|Имения у него было: семь тысяч мелкого скота, три тысячи верблюдов, пятьсот пар волов и пятьсот ослиц и весьма много прислуги; и был человек этот знаменитее всех сынов Востока.
JOB|1|4|Сыновья его сходились, делая пиры каждый в своем доме в свой день, и посылали и приглашали трех сестер своих есть и пить с ними.
JOB|1|5|Когда круг пиршественных дней совершался, Иов посылал [за ними] и освящал их и, вставая рано утром, возносил всесожжения по числу всех их. Ибо говорил Иов: может быть, сыновья мои согрешили и похулили Бога в сердце своем. Так делал Иов во все [такие] дни.
JOB|1|6|И был день, когда пришли сыны Божии предстать пред Господа; между ними пришел и сатана.
JOB|1|7|И сказал Господь сатане: откуда ты пришел? И отвечал сатана Господу и сказал: я ходил по земле и обошел ее.
JOB|1|8|И сказал Господь сатане: обратил ли ты внимание твое на раба Моего Иова? ибо нет такого, как он, на земле: человек непорочный, справедливый, богобоязненный и удаляющийся от зла.
JOB|1|9|И отвечал сатана Господу и сказал: разве даром богобоязнен Иов?
JOB|1|10|Не Ты ли кругом оградил его и дом его и все, что у него? Дело рук его Ты благословил, и стада его распространяются по земле;
JOB|1|11|но простри руку Твою и коснись всего, что у него, – благословит ли он Тебя?
JOB|1|12|И сказал Господь сатане: вот, все, что у него, в руке твоей; только на него не простирай руки твоей. И отошел сатана от лица Господня.
JOB|1|13|И был день, когда сыновья его и дочери его ели и вино пили в доме первородного брата своего.
JOB|1|14|И [вот], приходит вестник к Иову и говорит:
JOB|1|15|волы орали, и ослицы паслись подле них, как напали Савеяне и взяли их, а отроков поразили острием меча; и спасся только я один, чтобы возвестить тебе.
JOB|1|16|Еще он говорил, как приходит другой и сказывает: огонь Божий упал с неба и опалил овец и отроков и пожрал их; и спасся только я один, чтобы возвестить тебе.
JOB|1|17|Еще он говорил, как приходит другой и сказывает: Халдеи расположились тремя отрядами и бросились на верблюдов и взяли их, а отроков поразили острием меча; и спасся только я один, чтобы возвестить тебе.
JOB|1|18|Еще этот говорил, приходит другой и сказывает: сыновья твои и дочери твои ели и вино пили в доме первородного брата своего;
JOB|1|19|и вот, большой ветер пришел от пустыни и охватил четыре угла дома, и дом упал на отроков, и они умерли; и спасся только я один, чтобы возвестить тебе.
JOB|1|20|Тогда Иов встал и разодрал верхнюю одежду свою, остриг голову свою и пал на землю и поклонился
JOB|1|21|и сказал: наг я вышел из чрева матери моей, наг и возвращусь. Господь дал, Господь и взял; да будет имя Господне благословенно!
JOB|1|22|Во всем этом не согрешил Иов и не произнес ничего неразумного о Боге.
JOB|2|1|Был день, когда пришли сыны Божии предстать пред Господа; между ними пришел и сатана предстать пред Господа.
JOB|2|2|И сказал Господь сатане: откуда ты пришел? И отвечал сатана Господу и сказал: я ходил по земле и обошел ее.
JOB|2|3|И сказал Господь сатане: обратил ли ты внимание твое на раба Моего Иова? ибо нет такого, как он, на земле: человек непорочный, справедливый, богобоязненный и удаляющийся от зла, и доселе тверд в своей непорочности; а ты возбуждал Меня против него, чтобы погубить его безвинно.
JOB|2|4|И отвечал сатана Господу и сказал: кожу за кожу, а за жизнь свою отдаст человек все, что есть у него;
JOB|2|5|но простри руку Твою и коснись кости его и плоти его, – благословит ли он Тебя?
JOB|2|6|И сказал Господь сатане: вот, он в руке твоей, только душу его сбереги.
JOB|2|7|И отошел сатана от лица Господня и поразил Иова проказою лютою от подошвы ноги его по самое темя его.
JOB|2|8|И взял он себе черепицу, чтобы скоблить себя ею, и сел в пепел.
JOB|2|9|И сказала ему жена его: ты все еще тверд в непорочности твоей! похули Бога и умри.
JOB|2|10|Но он сказал ей: ты говоришь как одна из безумных: неужели доброе мы будем принимать от Бога, а злого не будем принимать? Во всем этом не согрешил Иов устами своими.
JOB|2|11|И услышали трое друзей Иова о всех этих несчастьях, постигших его, и пошли каждый из своего места: Елифаз Феманитянин, Вилдад Савхеянин и Софар Наамитянин, и сошлись, чтобы идти вместе сетовать с ним и утешать его.
JOB|2|12|И подняв глаза свои издали, они не узнали его; и возвысили голос свой и зарыдали; и разодрал каждый верхнюю одежду свою, и бросали пыль над головами своими к небу.
JOB|2|13|И сидели с ним на земле семь дней и семь ночей; и никто не говорил ему ни слова, ибо видели, что страдание его весьма велико.
JOB|3|1|После того открыл Иов уста свои и проклял день свой.
JOB|3|2|И начал Иов и сказал:
JOB|3|3|погибни день, в который я родился, и ночь, в которую сказано: зачался человек!
JOB|3|4|День тот да будет тьмою; да не взыщет его Бог свыше, и да не воссияет над ним свет!
JOB|3|5|Да омрачит его тьма и тень смертная, да обложит его туча, да страшатся его, как палящего зноя!
JOB|3|6|Ночь та, – да обладает ею мрак, да не сочтется она в днях года, да не войдет в число месяцев!
JOB|3|7|О! ночь та – да будет она безлюдна; да не войдет в нее веселье!
JOB|3|8|Да проклянут ее проклинающие день, способные разбудить левиафана!
JOB|3|9|Да померкнут звезды рассвета ее: пусть ждет она света, и он не приходит, и да не увидит она ресниц денницы
JOB|3|10|за то, что не затворила дверей чрева [матери] моей и не сокрыла горести от очей моих!
JOB|3|11|Для чего не умер я, выходя из утробы, и не скончался, когда вышел из чрева?
JOB|3|12|Зачем приняли меня колени? зачем было мне сосать сосцы?
JOB|3|13|Теперь бы лежал я и почивал; спал бы, и мне было бы покойно
JOB|3|14|с царями и советниками земли, которые застраивали для себя пустыни,
JOB|3|15|или с князьями, у которых было золото, и которые наполняли домы свои серебром;
JOB|3|16|или, как выкидыш сокрытый, я не существовал бы, как младенцы, не увидевшие света.
JOB|3|17|Там беззаконные перестают наводить страх, и там отдыхают истощившиеся в силах.
JOB|3|18|Там узники вместе наслаждаются покоем и не слышат криков приставника.
JOB|3|19|Малый и великий там равны, и раб свободен от господина своего.
JOB|3|20|На что дан страдальцу свет, и жизнь огорченным душею,
JOB|3|21|которые ждут смерти, и нет ее, которые вырыли бы ее охотнее, нежели клад,
JOB|3|22|обрадовались бы до восторга, восхитились бы, что нашли гроб?
JOB|3|23|[На что дан свет] человеку, которого путь закрыт, и которого Бог окружил мраком?
JOB|3|24|Вздохи мои предупреждают хлеб мой, и стоны мои льются, как вода,
JOB|3|25|ибо ужасное, чего я ужасался, то и постигло меня; и чего я боялся, то и пришло ко мне.
JOB|3|26|Нет мне мира, нет покоя, нет отрады: постигло несчастье.
JOB|4|1|И отвечал Елифаз Феманитянин и сказал:
JOB|4|2|[если] попытаемся мы [сказать] к тебе слово, – не тяжело ли будет тебе? Впрочем кто может возбранить слову!
JOB|4|3|Вот, ты наставлял многих и опустившиеся руки поддерживал,
JOB|4|4|падающего восставляли слова твои, и гнущиеся колени ты укреплял.
JOB|4|5|А теперь дошло до тебя, и ты изнемог; коснулось тебя, и ты упал духом.
JOB|4|6|Богобоязненность твоя не должна ли быть твоею надеждою, и непорочность путей твоих – упованием твоим?
JOB|4|7|Вспомни же, погибал ли кто невинный, и где праведные бывали искореняемы?
JOB|4|8|Как я видал, то оравшие нечестие и сеявшие зло пожинают его;
JOB|4|9|от дуновения Божия погибают и от духа гнева Его исчезают.
JOB|4|10|Рев льва и голос рыкающего [умолкает], и зубы скимнов сокрушаются;
JOB|4|11|могучий лев погибает без добычи, и дети львицы рассеиваются.
JOB|4|12|И вот, ко мне тайно принеслось слово, и ухо мое приняло нечто от него.
JOB|4|13|Среди размышлений о ночных видениях, когда сон находит на людей,
JOB|4|14|объял меня ужас и трепет и потряс все кости мои.
JOB|4|15|И дух прошел надо мною; дыбом стали волосы на мне.
JOB|4|16|Он стал, – но я не распознал вида его, – только облик был пред глазами моими; тихое веяние, – и я слышу голос:
JOB|4|17|человек праведнее ли Бога? и муж чище ли Творца своего?
JOB|4|18|Вот, Он и слугам Своим не доверяет и в Ангелах Своих усматривает недостатки:
JOB|4|19|тем более – в обитающих в храминах из брения, которых основание прах, которые истребляются скорее моли.
JOB|4|20|Между утром и вечером они распадаются; не увидишь, как они вовсе исчезнут.
JOB|4|21|Не погибают ли с ними и достоинства их? Они умирают, не достигнув мудрости.
JOB|5|1|Взывай, если есть отвечающий тебе. И к кому из святых обратишься ты?
JOB|5|2|Так, глупца убивает гневливость, и несмысленного губит раздражительность.
JOB|5|3|Видел я, как глупец укореняется, и тотчас проклял дом его.
JOB|5|4|Дети его далеки от счастья, их будут бить у ворот, и не будет заступника.
JOB|5|5|Жатву его съест голодный и из–за терна возьмет ее, и жаждущие поглотят имущество его.
JOB|5|6|Так, не из праха выходит горе, и не из земли вырастает беда;
JOB|5|7|но человек рождается на страдание, [как] искры, чтобы устремляться вверх.
JOB|5|8|Но я к Богу обратился бы, предал бы дело мое Богу,
JOB|5|9|Который творит дела великие и неисследимые, чудные без числа,
JOB|5|10|дает дождь на лице земли и посылает воды на лице полей;
JOB|5|11|униженных поставляет на высоту, и сетующие возносятся во спасение.
JOB|5|12|Он разрушает замыслы коварных, и руки их не довершают предприятия.
JOB|5|13|Он уловляет мудрецов их же лукавством, и совет хитрых становится тщетным:
JOB|5|14|днем они встречают тьму и в полдень ходят ощупью, как ночью.
JOB|5|15|Он спасает бедного от меча, от уст их и от руки сильного.
JOB|5|16|И есть несчастному надежда, и неправда затворяет уста свои.
JOB|5|17|Блажен человек, которого вразумляет Бог, и потому наказания Вседержителева не отвергай,
JOB|5|18|ибо Он причиняет раны и Сам обвязывает их; Он поражает, и Его же руки врачуют.
JOB|5|19|В шести бедах спасет тебя, и в седьмой не коснется тебя зло.
JOB|5|20|Во время голода избавит тебя от смерти, и на войне – от руки меча.
JOB|5|21|От бича языка укроешь себя и не убоишься опустошения, когда оно придет.
JOB|5|22|Опустошению и голоду посмеешься и зверей земли не убоишься,
JOB|5|23|ибо с камнями полевыми у тебя союз, и звери полевые в мире с тобою.
JOB|5|24|И узнаешь, что шатер твой в безопасности, и будешь смотреть за домом твоим, и не согрешишь.
JOB|5|25|И увидишь, что семя твое многочисленно, и отрасли твои, как трава на земле.
JOB|5|26|Войдешь во гроб в зрелости, как укладываются снопы пшеницы в свое время.
JOB|5|27|Вот, что мы дознали; так оно и есть: выслушай это и заметь для себя.
JOB|6|1|И отвечал Иов и сказал:
JOB|6|2|о, если бы верно взвешены были вопли мои, и вместе с ними положили на весы страдание мое!
JOB|6|3|Оно верно перетянуло бы песок морей! От того слова мои неистовы.
JOB|6|4|Ибо стрелы Вседержителя во мне; яд их пьет дух мой; ужасы Божии ополчились против меня.
JOB|6|5|Ревет ли дикий осел на траве? мычит ли бык у месива своего?
JOB|6|6|Едят ли безвкусное без соли, и есть ли вкус в яичном белке?
JOB|6|7|До чего не хотела коснуться душа моя, то составляет отвратительную пищу мою.
JOB|6|8|О, когда бы сбылось желание мое и чаяние мое исполнил Бог!
JOB|6|9|О, если бы благоволил Бог сокрушить меня, простер руку Свою и сразил меня!
JOB|6|10|Это было бы еще отрадою мне, и я крепился бы в моей беспощадной болезни, ибо я не отвергся изречений Святаго.
JOB|6|11|Что за сила у меня, чтобы надеяться мне? и какой конец, чтобы длить мне жизнь мою?
JOB|6|12|Твердость ли камней твердость моя? и медь ли плоть моя?
JOB|6|13|Есть ли во мне помощь для меня, и есть ли для меня какая опора?
JOB|6|14|К страждущему должно быть сожаление от друга его, если только он не оставил страха к Вседержителю.
JOB|6|15|Но братья мои неверны, как поток, как быстро текущие ручьи,
JOB|6|16|которые черны от льда и в которых скрывается снег.
JOB|6|17|Когда становится тепло, они умаляются, а во время жары исчезают с мест своих.
JOB|6|18|Уклоняют они направление путей своих, заходят в пустыню и теряются;
JOB|6|19|смотрят на них дороги Фемайские, надеются на них пути Савейские,
JOB|6|20|но остаются пристыженными в своей надежде; приходят туда и от стыда краснеют.
JOB|6|21|Так и вы теперь ничто: увидели страшное и испугались.
JOB|6|22|Говорил ли я: дайте мне, или от достатка вашего заплатите за меня;
JOB|6|23|и избавьте меня от руки врага, и от руки мучителей выкупите меня?
JOB|6|24|Научите меня, и я замолчу; укажите, в чем я погрешил.
JOB|6|25|Как сильны слова правды! Но что доказывают обличения ваши?
JOB|6|26|Вы придумываете речи для обличения? На ветер пускаете слова ваши.
JOB|6|27|Вы нападаете на сироту и роете яму другу вашему.
JOB|6|28|Но прошу вас, взгляните на меня; буду ли я говорить ложь пред лицем вашим?
JOB|6|29|Пересмотрите, есть ли неправда? пересмотрите, – правда моя.
JOB|6|30|Есть ли на языке моем неправда? Неужели гортань моя не может различить горечи?
JOB|7|1|Не определено ли человеку время на земле, и дни его не то же ли, что дни наемника?
JOB|7|2|Как раб жаждет тени, и как наемник ждет окончания работы своей,
JOB|7|3|так я получил в удел месяцы суетные, и ночи горестные отчислены мне.
JOB|7|4|Когда ложусь, то говорю: "когда–то встану?", а вечер длится, и я ворочаюсь досыта до самого рассвета.
JOB|7|5|Тело мое одето червями и пыльными струпами; кожа моя лопается и гноится.
JOB|7|6|Дни мои бегут скорее челнока и кончаются без надежды.
JOB|7|7|Вспомни, что жизнь моя дуновение, что око мое не возвратится видеть доброе.
JOB|7|8|Не увидит меня око видевшего меня; очи Твои на меня, – и нет меня.
JOB|7|9|Редеет облако и уходит; так нисшедший в преисподнюю не выйдет,
JOB|7|10|не возвратится более в дом свой, и место его не будет уже знать его.
JOB|7|11|Не буду же я удерживать уст моих; буду говорить в стеснении духа моего; буду жаловаться в горести души моей.
JOB|7|12|Разве я море или морское чудовище, что Ты поставил надо мною стражу?
JOB|7|13|Когда подумаю: утешит меня постель моя, унесет горесть мою ложе мое,
JOB|7|14|ты страшишь меня снами и видениями пугаешь меня;
JOB|7|15|и душа моя желает лучше прекращения дыхания, лучше смерти, нежели [сбережения] костей моих.
JOB|7|16|Опротивела мне жизнь. Не вечно жить мне. Отступи от меня, ибо дни мои суета.
JOB|7|17|Что такое человек, что Ты столько ценишь его и обращаешь на него внимание Твое,
JOB|7|18|посещаешь его каждое утро, каждое мгновение испытываешь его?
JOB|7|19|Доколе же Ты не оставишь, доколе не отойдешь от меня, доколе не дашь мне проглотить слюну мою?
JOB|7|20|Если я согрешил, то что я сделаю Тебе, страж человеков! Зачем Ты поставил меня противником Себе, так что я стал самому себе в тягость?
JOB|7|21|И зачем бы не простить мне греха и не снять с меня беззакония моего? ибо, вот, я лягу в прахе; завтра поищешь меня, и меня нет.
JOB|8|1|И отвечал Вилдад Савхеянин и сказал:
JOB|8|2|долго ли ты будешь говорить так? – слова уст твоих бурный ветер!
JOB|8|3|Неужели Бог извращает суд, и Вседержитель превращает правду?
JOB|8|4|Если сыновья твои согрешили пред Ним, то Он и предал их в руку беззакония их.
JOB|8|5|Если же ты взыщешь Бога и помолишься Вседержителю,
JOB|8|6|и если ты чист и прав, то Он ныне же встанет над тобою и умиротворит жилище правды твоей.
JOB|8|7|И если вначале у тебя было мало, то впоследствии будет весьма много.
JOB|8|8|Ибо спроси у прежних родов и вникни в наблюдения отцов их;
JOB|8|9|а мы – вчерашние и ничего не знаем, потому что наши дни на земле тень.
JOB|8|10|Вот они научат тебя, скажут тебе и от сердца своего произнесут слова:
JOB|8|11|поднимается ли тростник без влаги? растет ли камыш без воды?
JOB|8|12|Еще он в свежести своей и не срезан, а прежде всякой травы засыхает.
JOB|8|13|Таковы пути всех забывающих Бога, и надежда лицемера погибнет;
JOB|8|14|упование его подсечено, и уверенность его – дом паука.
JOB|8|15|Обопрется о дом свой и не устоит; ухватится за него и не удержится.
JOB|8|16|Зеленеет он пред солнцем, за сад простираются ветви его;
JOB|8|17|в кучу [камней] вплетаются корни его, между камнями врезываются.
JOB|8|18|Но когда вырвут его с места его, оно откажется от него: "я не видало тебя!"
JOB|8|19|Вот радость пути его! а из земли вырастают другие.
JOB|8|20|Видишь, Бог не отвергает непорочного и не поддерживает руки злодеев.
JOB|8|21|Он еще наполнит смехом уста твои и губы твои радостным восклицанием.
JOB|8|22|Ненавидящие тебя облекутся в стыд, и шатра нечестивых не станет.
JOB|9|1|И отвечал Иов и сказал:
JOB|9|2|правда! знаю, что так; но как оправдается человек пред Богом?
JOB|9|3|Если захочет вступить в прение с Ним, то не ответит Ему ни на одно из тысячи.
JOB|9|4|Премудр сердцем и могущ силою; кто восставал против Него и оставался в покое?
JOB|9|5|Он передвигает горы, и не узнают их: Он превращает их в гневе Своем;
JOB|9|6|сдвигает землю с места ее, и столбы ее дрожат;
JOB|9|7|скажет солнцу, – и не взойдет, и на звезды налагает печать.
JOB|9|8|Он один распростирает небеса и ходит по высотам моря;
JOB|9|9|сотворил Ас, Кесиль и Хима и тайники юга;
JOB|9|10|делает великое, неисследимое и чудное без числа!
JOB|9|11|Вот, Он пройдет предо мною, и не увижу Его; пронесется и не замечу Его.
JOB|9|12|Возьмет, и кто возбранит Ему? кто скажет Ему: что Ты делаешь?
JOB|9|13|Бог не отвратит гнева Своего; пред Ним падут поборники гордыни.
JOB|9|14|Тем более могу ли я отвечать Ему и приискивать себе слова пред Ним?
JOB|9|15|Хотя бы я и прав был, но не буду отвечать, а буду умолять Судию моего.
JOB|9|16|Если бы я воззвал, и Он ответил мне, – я не поверил бы, что голос мой услышал Тот,
JOB|9|17|Кто в вихре разит меня и умножает безвинно мои раны,
JOB|9|18|не дает мне перевести духа, но пресыщает меня горестями.
JOB|9|19|Если [действовать] силою, то Он могуществен; если судом, кто сведет меня с Ним?
JOB|9|20|Если я буду оправдываться, то мои же уста обвинят меня; [если] я невинен, то Он признает меня виновным.
JOB|9|21|Невинен я; не хочу знать души моей, презираю жизнь мою.
JOB|9|22|Все одно; поэтому я сказал, что Он губит и непорочного и виновного.
JOB|9|23|Если этого поражает Он бичом вдруг, то пытке невинных посмевается.
JOB|9|24|Земля отдана в руки нечестивых; лица судей ее Он закрывает. Если не Он, то кто же?
JOB|9|25|Дни мои быстрее гонца, – бегут, не видят добра,
JOB|9|26|несутся, как легкие ладьи, как орел стремится на добычу.
JOB|9|27|Если сказать мне: забуду я жалобы мои, отложу мрачный вид свой и ободрюсь;
JOB|9|28|то трепещу всех страданий моих, зная, что Ты не объявишь меня невинным.
JOB|9|29|Если же я виновен, то для чего напрасно томлюсь?
JOB|9|30|Хотя бы я омылся и снежною водою и совершенно очистил руки мои,
JOB|9|31|то и тогда Ты погрузишь меня в грязь, и возгнушаются мною одежды мои.
JOB|9|32|Ибо Он не человек, как я, чтоб я мог отвечать Ему и идти вместе с Ним на суд!
JOB|9|33|Нет между нами посредника, который положил бы руку свою на обоих нас.
JOB|9|34|Да отстранит Он от меня жезл Свой, и страх Его да не ужасает меня, –
JOB|9|35|и тогда я буду говорить и не убоюсь Его, ибо я не таков сам в себе.
JOB|10|1|Опротивела душе моей жизнь моя; предамся печали моей; буду говорить в горести души моей.
JOB|10|2|Скажу Богу: не обвиняй меня; объяви мне, за что Ты со мною борешься?
JOB|10|3|Хорошо ли для Тебя, что Ты угнетаешь, что презираешь дело рук Твоих, а на совет нечестивых посылаешь свет?
JOB|10|4|Разве у Тебя плотские очи, и Ты смотришь, как смотрит человек?
JOB|10|5|Разве дни Твои, как дни человека, или лета Твои, как дни мужа,
JOB|10|6|что Ты ищешь порока во мне и допытываешься греха во мне,
JOB|10|7|хотя знаешь, что я не беззаконник, и что некому избавить меня от руки Твоей?
JOB|10|8|Твои руки трудились надо мною и образовали всего меня кругом, – и Ты губишь меня?
JOB|10|9|Вспомни, что Ты, как глину, обделал меня, и в прах обращаешь меня?
JOB|10|10|Не Ты ли вылил меня, как молоко, и, как творог, сгустил меня,
JOB|10|11|кожею и плотью одел меня, костями и жилами скрепил меня,
JOB|10|12|жизнь и милость даровал мне, и попечение Твое хранило дух мой?
JOB|10|13|Но и то скрывал Ты в сердце Своем, – знаю, что это было у Тебя, –
JOB|10|14|что если я согрешу, Ты заметишь и не оставишь греха моего без наказания.
JOB|10|15|Если я виновен, горе мне! если и прав, то не осмелюсь поднять головы моей. Я пресыщен унижением; взгляни на бедствие мое:
JOB|10|16|оно увеличивается. Ты гонишься за мною, как лев, и снова нападаешь на меня и чудным являешься во мне.
JOB|10|17|Выводишь новых свидетелей Твоих против меня; усиливаешь гнев Твой на меня; и беды, одни за другими, ополчаются против меня.
JOB|10|18|И зачем Ты вывел меня из чрева? пусть бы я умер, когда еще ничей глаз не видел меня;
JOB|10|19|пусть бы я, как небывший, из чрева перенесен был во гроб!
JOB|10|20|Не малы ли дни мои? Оставь, отступи от меня, чтобы я немного ободрился,
JOB|10|21|прежде нежели отойду, – и уже не возвращусь, – в страну тьмы и сени смертной,
JOB|10|22|в страну мрака, каков есть мрак тени смертной, где нет устройства, [где] темно, как самая тьма.
JOB|11|1|И отвечал Софар Наамитянин и сказал:
JOB|11|2|разве на множество слов нельзя дать ответа, и разве человек многоречивый прав?
JOB|11|3|Пустословие твое заставит ли молчать мужей, чтобы ты глумился, и некому было постыдить тебя?
JOB|11|4|Ты сказал: суждение мое верно, и чист я в очах Твоих.
JOB|11|5|Но если бы Бог возглаголал и отверз уста Свои к тебе
JOB|11|6|и открыл тебе тайны премудрости, что тебе вдвое больше следовало бы понести! Итак знай, что Бог для тебя некоторые из беззаконий твоих предал забвению.
JOB|11|7|Можешь ли ты исследованием найти Бога? Можешь ли совершенно постигнуть Вседержителя?
JOB|11|8|Он превыше небес, – что можешь сделать? глубже преисподней, – что можешь узнать?
JOB|11|9|Длиннее земли мера Его и шире моря.
JOB|11|10|Если Он пройдет и заключит кого в оковы и представит на суд, то кто отклонит Его?
JOB|11|11|Ибо Он знает людей лживых и видит беззаконие, и оставит ли его без внимания?
JOB|11|12|Но пустой человек мудрствует, хотя человек рождается подобно дикому осленку.
JOB|11|13|Если ты управишь сердце твое и прострешь к Нему руки твои,
JOB|11|14|и если есть порок в руке твоей, а ты удалишь его и не дашь беззаконию обитать в шатрах твоих,
JOB|11|15|то поднимешь незапятнанное лице твое и будешь тверд и не будешь бояться.
JOB|11|16|Тогда забудешь горе: как о воде протекшей, будешь вспоминать о нем.
JOB|11|17|И яснее полдня пойдет жизнь твоя; просветлеешь, как утро.
JOB|11|18|И будешь спокоен, ибо есть надежда; ты огражден, и можешь спать безопасно.
JOB|11|19|Будешь лежать, и не будет устрашающего, и многие будут заискивать у тебя.
JOB|11|20|глаза беззаконных истают, и убежище пропадет у них, и надежда их исчезнет.
JOB|12|1|И отвечал Иов и сказал:
JOB|12|2|подлинно, [только] вы люди, и с вами умрет мудрость!
JOB|12|3|И у меня [есть] сердце, как у вас; не ниже я вас; и кто не знает того же?
JOB|12|4|Посмешищем стал я для друга своего, я, который взывал к Богу, и которому Он отвечал, посмешищем – [человек] праведный, непорочный.
JOB|12|5|Так презрен по мыслям сидящего в покое факел, приготовленный для спотыкающихся ногами.
JOB|12|6|Покойны шатры у грабителей и безопасны у раздражающих Бога, которые как бы Бога носят в руках своих.
JOB|12|7|И подлинно: спроси у скота, и научит тебя, у птицы небесной, и возвестит тебе;
JOB|12|8|или побеседуй с землею, и наставит тебя, и скажут тебе рыбы морские.
JOB|12|9|Кто во всем этом не узнает, что рука Господа сотворила сие?
JOB|12|10|В Его руке душа всего живущего и дух всякой человеческой плоти.
JOB|12|11|Не ухо ли разбирает слова, и не язык ли распознает вкус пищи?
JOB|12|12|В старцах – мудрость, и в долголетних – разум.
JOB|12|13|У Него премудрость и сила; Его совет и разум.
JOB|12|14|Что Он разрушит, то не построится; кого Он заключит, тот не высвободится.
JOB|12|15|Остановит воды, и все высохнет; пустит их, и превратят землю.
JOB|12|16|У Него могущество и премудрость, пред Ним заблуждающийся и вводящий в заблуждение.
JOB|12|17|Он приводит советников в необдуманность и судей делает глупыми.
JOB|12|18|Он лишает перевязей царей и поясом обвязывает чресла их;
JOB|12|19|князей лишает достоинства и низвергает храбрых;
JOB|12|20|отнимает язык у велеречивых и старцев лишает смысла;
JOB|12|21|покрывает стыдом знаменитых и силу могучих ослабляет;
JOB|12|22|открывает глубокое из среды тьмы и выводит на свет тень смертную;
JOB|12|23|умножает народы и истребляет их; рассевает народы и собирает их;
JOB|12|24|отнимает ум у глав народа земли и оставляет их блуждать в пустыне, где нет пути:
JOB|12|25|ощупью ходят они во тьме без света и шатаются, как пьяные.
JOB|13|1|Вот, все [это] видело око мое, слышало ухо мое и заметило для себя.
JOB|13|2|Сколько знаете вы, знаю и я: не ниже я вас.
JOB|13|3|Но я к Вседержителю хотел бы говорить и желал бы состязаться с Богом.
JOB|13|4|А вы сплетчики лжи; все вы бесполезные врачи.
JOB|13|5|О, если бы вы только молчали! это было бы [вменено] вам в мудрость.
JOB|13|6|Выслушайте же рассуждения мои и вникните в возражение уст моих.
JOB|13|7|Надлежало ли вам ради Бога говорить неправду и для Него говорить ложь?
JOB|13|8|Надлежало ли вам быть лицеприятными к Нему и за Бога так препираться?
JOB|13|9|Хорошо ли будет, когда Он испытает вас? Обманете ли Его, как обманывают человека?
JOB|13|10|Строго накажет Он вас, хотя вы и скрытно лицемерите.
JOB|13|11|Неужели величие Его не устрашает вас, и страх Его не нападает на вас?
JOB|13|12|Напоминания ваши подобны пеплу; оплоты ваши – оплоты глиняные.
JOB|13|13|Замолчите предо мною, и я буду говорить, что бы ни постигло меня.
JOB|13|14|Для чего мне терзать тело мое зубами моими и душу мою полагать в руку мою?
JOB|13|15|Вот, Он убивает меня, но я буду надеяться; я желал бы только отстоять пути мои пред лицем Его!
JOB|13|16|И это уже в оправдание мне, потому что лицемер не пойдет пред лице Его!
JOB|13|17|Выслушайте внимательно слово мое и объяснение мое ушами вашими.
JOB|13|18|Вот, я завел судебное дело: знаю, что буду прав.
JOB|13|19|Кто в состоянии оспорить меня? Ибо я скоро умолкну и испущу дух.
JOB|13|20|Двух только [вещей] не делай со мною, и тогда я не буду укрываться от лица Твоего:
JOB|13|21|удали от меня руку Твою, и ужас Твой да не потрясает меня.
JOB|13|22|Тогда зови, и я буду отвечать, или буду говорить я, а Ты отвечай мне.
JOB|13|23|Сколько у меня пороков и грехов? покажи мне беззаконие мое и грех мой.
JOB|13|24|Для чего скрываешь лице Твое и считаешь меня врагом Тебе?
JOB|13|25|Не сорванный ли листок Ты сокрушаешь и не сухую ли соломинку преследуешь?
JOB|13|26|Ибо Ты пишешь на меня горькое и вменяешь мне грехи юности моей,
JOB|13|27|и ставишь в колоду ноги мои и подстерегаешь все стези мои, – гонишься по следам ног моих.
JOB|13|28|А он, как гниль, распадается, как одежда, изъеденная молью.
JOB|14|1|Человек, рожденный женою, краткодневен и пресыщен печалями:
JOB|14|2|как цветок, он выходит и опадает; убегает, как тень, и не останавливается.
JOB|14|3|И на него–то Ты отверзаешь очи Твои, и меня ведешь на суд с Тобою?
JOB|14|4|Кто родится чистым от нечистого? Ни один.
JOB|14|5|Если дни ему определены, и число месяцев его у Тебя, если Ты положил ему предел, которого он не перейдет,
JOB|14|6|то уклонись от него: пусть он отдохнет, доколе не окончит, как наемник, дня своего.
JOB|14|7|Для дерева есть надежда, что оно, если и будет срублено, снова оживет, и отрасли от него [выходить] не перестанут:
JOB|14|8|если и устарел в земле корень его, и пень его замер в пыли,
JOB|14|9|но, лишь почуяло воду, оно дает отпрыски и пускает ветви, как бы вновь посаженное.
JOB|14|10|А человек умирает и распадается; отошел, и где он?
JOB|14|11|Уходят воды из озера, и река иссякает и высыхает:
JOB|14|12|так человек ляжет и не станет; до скончания неба он не пробудится и не воспрянет от сна своего.
JOB|14|13|О, если бы Ты в преисподней сокрыл меня и укрывал меня, пока пройдет гнев Твой, положил мне срок и потом вспомнил обо мне!
JOB|14|14|Когда умрет человек, то будет ли он опять жить? Во все дни определенного мне времени я ожидал бы, пока придет мне смена.
JOB|14|15|Воззвал бы Ты, и я дал бы Тебе ответ, и Ты явил бы благоволение творению рук Твоих;
JOB|14|16|ибо тогда Ты исчислял бы шаги мои и не подстерегал бы греха моего;
JOB|14|17|в свитке было бы запечатано беззаконие мое, и Ты закрыл бы вину мою.
JOB|14|18|Но гора падая разрушается, и скала сходит с места своего;
JOB|14|19|вода стирает камни; разлив ее смывает земную пыль: так и надежду человека Ты уничтожаешь.
JOB|14|20|Теснишь его до конца, и он уходит; изменяешь ему лице и отсылаешь его.
JOB|14|21|В чести ли дети его – он не знает, унижены ли – он не замечает;
JOB|14|22|но плоть его на нем болит, и душа его в нем страдает.
JOB|15|1|И отвечал Елифаз Феманитянин и сказал:
JOB|15|2|станет ли мудрый отвечать знанием пустым и наполнять чрево свое ветром палящим,
JOB|15|3|оправдываться словами бесполезными и речью, не имеющею никакой силы?
JOB|15|4|Да ты отложил и страх и за малость считаешь речь к Богу.
JOB|15|5|Нечестие твое настроило так уста твои, и ты избрал язык лукавых.
JOB|15|6|Тебя обвиняют уста твои, а не я, и твой язык говорит против тебя.
JOB|15|7|Разве ты первым человеком родился и прежде холмов создан?
JOB|15|8|Разве совет Божий ты слышал и привлек к себе премудрость?
JOB|15|9|Что знаешь ты, чего бы не знали мы? что разумеешь ты, чего не было бы и у нас?
JOB|15|10|И седовласый и старец есть между нами, днями превышающий отца твоего.
JOB|15|11|Разве малость для тебя утешения Божии? И это неизвестно тебе?
JOB|15|12|К чему порывает тебя сердце твое, и к чему так гордо смотришь?
JOB|15|13|Что устремляешь против Бога дух твой и устами твоими произносишь такие речи?
JOB|15|14|Что такое человек, чтоб быть ему чистым, и чтобы рожденному женщиною быть праведным?
JOB|15|15|Вот, Он и святым Своим не доверяет, и небеса нечисты в очах Его:
JOB|15|16|тем больше нечист и растлен человек, пьющий беззаконие, как воду.
JOB|15|17|Я буду говорить тебе, слушай меня; я расскажу тебе, что видел,
JOB|15|18|что слышали мудрые и не скрыли слышанного от отцов своих,
JOB|15|19|которым одним отдана была земля, и среди которых чужой не ходил.
JOB|15|20|Нечестивый мучит себя во все дни свои, и число лет закрыто от притеснителя;
JOB|15|21|звук ужасов в ушах его; среди мира идет на него губитель.
JOB|15|22|Он не надеется спастись от тьмы; видит пред собою меч.
JOB|15|23|Он скитается за куском хлеба повсюду; знает, что уже готов, в руках у него день тьмы.
JOB|15|24|Устрашает его нужда и теснота; одолевает его, как царь, приготовившийся к битве,
JOB|15|25|за то, что он простирал против Бога руку свою и противился Вседержителю,
JOB|15|26|устремлялся против Него с [гордою] выею, под толстыми щитами своими;
JOB|15|27|потому что он покрыл лице свое жиром своим и обложил туком лядвеи свои.
JOB|15|28|И он селится в городах разоренных, в домах, в которых не живут, которые обречены на развалины.
JOB|15|29|Не пребудет он богатым, и не уцелеет имущество его, и не распрострется по земле приобретение его.
JOB|15|30|Не уйдет от тьмы; отрасли его иссушит пламя и дуновением уст своих увлечет его.
JOB|15|31|Пусть не доверяет суете заблудший, ибо суета будет и воздаянием ему.
JOB|15|32|Не в свой день он скончается, и ветви его не будут зеленеть.
JOB|15|33|Сбросит он, как виноградная лоза, недозрелую ягоду свою и, как маслина, стряхнет цвет свой.
JOB|15|34|Так опустеет дом нечестивого, и огонь пожрет шатры мздоимства.
JOB|15|35|Он зачал зло и родил ложь, и утроба его приготовляет обман.
JOB|16|1|И отвечал Иов и сказал:
JOB|16|2|слышал я много такого; жалкие утешители все вы!
JOB|16|3|Будет ли конец ветреным словам? и что побудило тебя так отвечать?
JOB|16|4|И я мог бы так же говорить, как вы, если бы душа ваша была на месте души моей; ополчался бы на вас словами и кивал бы на вас головою моею;
JOB|16|5|подкреплял бы вас языком моим и движением губ утешал бы.
JOB|16|6|Говорю ли я, не утоляется скорбь моя; перестаю ли, что отходит от меня?
JOB|16|7|Но ныне Он изнурил меня. Ты разрушил всю семью мою.
JOB|16|8|Ты покрыл меня морщинами во свидетельство против меня; восстает на меня изможденность моя, в лицо укоряет меня.
JOB|16|9|Гнев Его терзает и враждует против меня, скрежещет на меня зубами своими; неприятель мой острит на меня глаза свои.
JOB|16|10|Разинули на меня пасть свою; ругаясь бьют меня по щекам; все сговорились против меня.
JOB|16|11|Предал меня Бог беззаконнику и в руки нечестивым бросил меня.
JOB|16|12|Я был спокоен, но Он потряс меня; взял меня за шею и избил меня и поставил меня целью для Себя.
JOB|16|13|Окружили меня стрельцы Его; Он рассекает внутренности мои и не щадит, пролил на землю желчь мою,
JOB|16|14|пробивает во мне пролом за проломом, бежит на меня, как ратоборец.
JOB|16|15|Вретище сшил я на кожу мою и в прах положил голову мою.
JOB|16|16|Лицо мое побагровело от плача, и на веждах моих тень смерти,
JOB|16|17|при всем том, что нет хищения в руках моих, и молитва моя чиста.
JOB|16|18|Земля! не закрой моей крови, и да не будет места воплю моему.
JOB|16|19|И ныне вот на небесах Свидетель мой, и Заступник мой в вышних!
JOB|16|20|Многоречивые друзья мои! К Богу слезит око мое.
JOB|16|21|О, если бы человек мог иметь состязание с Богом, как сын человеческий с ближним своим!
JOB|16|22|Ибо летам моим приходит конец, и я отхожу в путь невозвратный.
JOB|17|1|Дыхание мое ослабело; дни мои угасают; гробы предо мною.
JOB|17|2|Если бы не насмешки их, то и среди споров их око мое пребывало бы спокойно.
JOB|17|3|Заступись, поручись [Сам] за меня пред Собою! иначе кто поручится за меня?
JOB|17|4|Ибо Ты закрыл сердце их от разумения, и потому не дашь восторжествовать [им].
JOB|17|5|Кто обрекает друзей своих в добычу, у детей того глаза истают.
JOB|17|6|Он поставил меня притчею для народа и посмешищем для него.
JOB|17|7|Помутилось от горести око мое, и все члены мои, как тень.
JOB|17|8|Изумятся о сем праведные, и невинный вознегодует на лицемера.
JOB|17|9|Но праведник будет крепко держаться пути своего, и чистый руками будет больше и больше утверждаться.
JOB|17|10|Выслушайте, все вы, и подойдите; не найду я мудрого между вами.
JOB|17|11|Дни мои прошли; думы мои – достояние сердца моего – разбиты.
JOB|17|12|А они ночь [хотят] превратить в день, свет приблизить к лицу тьмы.
JOB|17|13|Если бы я и ожидать стал, то преисподняя – дом мой; во тьме постелю я постель мою;
JOB|17|14|гробу скажу: ты отец мой, червю: ты мать моя и сестра моя.
JOB|17|15|Где же после этого надежда моя? и ожидаемое мною кто увидит?
JOB|17|16|В преисподнюю сойдет она и будет покоиться со мною в прахе.
JOB|18|1|И отвечал Вилдад Савхеянин и сказал:
JOB|18|2|когда же положите вы конец таким речам? обдумайте, и потом будем говорить.
JOB|18|3|Зачем считаться нам за животных и быть униженными в собственных глазах ваших?
JOB|18|4|[О ты], раздирающий душу твою в гневе твоем! Неужели для тебя опустеть земле, и скале сдвинуться с места своего?
JOB|18|5|Да, свет у беззаконного потухнет, и не останется искры от огня его.
JOB|18|6|Померкнет свет в шатре его, и светильник его угаснет над ним.
JOB|18|7|Сократятся шаги могущества его, и низложит его собственный замысл его,
JOB|18|8|ибо он попадет в сеть своими ногами и по тенетам ходить будет.
JOB|18|9|Петля зацепит за ногу его, и грабитель уловит его.
JOB|18|10|Скрытно разложены по земле силки для него и западни на дороге.
JOB|18|11|Со всех сторон будут страшить его ужасы и заставят его бросаться туда и сюда.
JOB|18|12|Истощится от голода сила его, и гибель готова, сбоку у него.
JOB|18|13|Съест члены тела его, съест члены его первенец смерти.
JOB|18|14|Изгнана будет из шатра его надежда его, и это низведет его к царю ужасов.
JOB|18|15|Поселятся в шатре его, потому что он уже не его; жилище его посыпано будет серою.
JOB|18|16|Снизу подсохнут корни его, и сверху увянут ветви его.
JOB|18|17|Память о нем исчезнет с земли, и имени его не будет на площади.
JOB|18|18|Изгонят его из света во тьму и сотрут его с лица земли.
JOB|18|19|Ни сына его, ни внука не будет в народе его, и никого не останется в жилищах его.
JOB|18|20|О дне его ужаснутся потомки, и современники будут объяты трепетом.
JOB|18|21|Таковы жилища беззаконного, и таково место того, кто не знает Бога.
JOB|19|1|И отвечал Иов и сказал:
JOB|19|2|доколе будете мучить душу мою и терзать меня речами?
JOB|19|3|Вот, уже раз десять вы срамили меня и не стыдитесь теснить меня.
JOB|19|4|Если я и действительно погрешил, то погрешность моя при мне остается.
JOB|19|5|Если же вы хотите повеличаться надо мною и упрекнуть меня позором моим,
JOB|19|6|то знайте, что Бог ниспроверг меня и обложил меня Своею сетью.
JOB|19|7|Вот, я кричу: обида! и никто не слушает; вопию, и нет суда.
JOB|19|8|Он преградил мне дорогу, и не могу пройти, и на стези мои положил тьму.
JOB|19|9|Совлек с меня славу мою и снял венец с головы моей.
JOB|19|10|Кругом разорил меня, и я отхожу; и, как дерево, Он исторг надежду мою.
JOB|19|11|Воспылал на меня гневом Своим и считает меня между врагами Своими.
JOB|19|12|Полки Его пришли вместе и направили путь свой ко мне и расположились вокруг шатра моего.
JOB|19|13|Братьев моих Он удалил от меня, и знающие меня чуждаются меня.
JOB|19|14|Покинули меня близкие мои, и знакомые мои забыли меня.
JOB|19|15|Пришлые в доме моем и служанки мои чужим считают меня; посторонним стал я в глазах их.
JOB|19|16|Зову слугу моего, и он не откликается; устами моими я должен умолять его.
JOB|19|17|Дыхание мое опротивело жене моей, и я должен умолять ее ради детей чрева моего.
JOB|19|18|Даже малые дети презирают меня: поднимаюсь, и они издеваются надо мною.
JOB|19|19|Гнушаются мною все наперсники мои, и те, которых я любил, обратились против меня.
JOB|19|20|Кости мои прилипли к коже моей и плоти моей, и я остался только с кожею около зубов моих.
JOB|19|21|Помилуйте меня, помилуйте меня вы, друзья мои, ибо рука Божия коснулась меня.
JOB|19|22|Зачем и вы преследуете меня, как Бог, и плотью моею не можете насытиться?
JOB|19|23|О, если бы записаны были слова мои! Если бы начертаны были они в книге
JOB|19|24|резцом железным с оловом, – на вечное время на камне вырезаны были!
JOB|19|25|А я знаю, Искупитель мой жив, и Он в последний день восставит из праха распадающуюся кожу мою сию,
JOB|19|26|и я во плоти моей узрю Бога.
JOB|19|27|Я узрю Его сам; мои глаза, не глаза другого, увидят Его. Истаевает сердце мое в груди моей!
JOB|19|28|Вам надлежало бы сказать: зачем мы преследуем его? Как будто корень зла найден во мне.
JOB|19|29|Убойтесь меча, ибо меч есть отмститель неправды, и знайте, что есть суд.
JOB|20|1|И отвечал Софар Наамитянин и сказал:
JOB|20|2|размышления мои побуждают меня отвечать, и я поспешаю выразить их.
JOB|20|3|Упрек, позорный для меня, выслушал я, и дух разумения моего ответит за меня.
JOB|20|4|Разве не знаешь ты, что от века, – с того времени, как поставлен человек на земле, –
JOB|20|5|веселье беззаконных кратковременно, и радость лицемера мгновенна?
JOB|20|6|Хотя бы возросло до небес величие его, и голова его касалась облаков, –
JOB|20|7|как помет его, на веки пропадает он; видевшие его скажут: где он?
JOB|20|8|Как сон, улетит, и не найдут его; и, как ночное видение, исчезнет.
JOB|20|9|Глаз, видевший его, больше не увидит его, и уже не усмотрит его место его.
JOB|20|10|Сыновья его будут заискивать у нищих, и руки его возвратят похищенное им.
JOB|20|11|Кости его наполнены грехами юности его, и с ним лягут они в прах.
JOB|20|12|Если сладко во рту его зло, и он таит его под языком своим,
JOB|20|13|бережет и не бросает его, а держит его в устах своих,
JOB|20|14|то эта пища его в утробе его превратится в желчь аспидов внутри его.
JOB|20|15|Имение, которое он глотал, изблюет: Бог исторгнет его из чрева его.
JOB|20|16|Змеиный яд он сосет; умертвит его язык ехидны.
JOB|20|17|Не видать ему ручьев, рек, текущих медом и молоком!
JOB|20|18|Нажитое трудом возвратит, не проглотит; по мере имения его будет и расплата его, а он не порадуется.
JOB|20|19|Ибо он угнетал, отсылал бедных; захватывал домы, которых не строил;
JOB|20|20|не знал сытости во чреве своем и в жадности своей не щадил ничего.
JOB|20|21|Ничего не спаслось от обжорства его, зато не устоит счастье его.
JOB|20|22|В полноте изобилия будет тесно ему; всякая рука обиженного поднимется на него.
JOB|20|23|Когда будет чем наполнить утробу его, Он пошлет на него ярость гнева Своего и одождит на него болезни в плоти его.
JOB|20|24|Убежит ли он от оружия железного, – пронзит его лук медный;
JOB|20|25|станет вынимать [стрелу], – и она выйдет из тела, выйдет, сверкая сквозь желчь его; ужасы смерти найдут на него!
JOB|20|26|Все мрачное сокрыто внутри его; будет пожирать его огонь, никем не раздуваемый; зло постигнет и оставшееся в шатре его.
JOB|20|27|Небо откроет беззаконие его, и земля восстанет против него.
JOB|20|28|Исчезнет стяжание дома его; все расплывется в день гнева Его.
JOB|20|29|Вот удел человеку беззаконному от Бога и наследие, определенное ему Вседержителем!
JOB|21|1|И отвечал Иов и сказал:
JOB|21|2|выслушайте внимательно речь мою, и это будет мне утешением от вас.
JOB|21|3|Потерпите меня, и я буду говорить; а после того, как поговорю, насмехайся.
JOB|21|4|Разве к человеку речь моя? как же мне и не малодушествовать?
JOB|21|5|Посмотрите на меня и ужаснитесь, и положите перст на уста.
JOB|21|6|Лишь только я вспомню, – содрогаюсь, и трепет объемлет тело мое.
JOB|21|7|Почему беззаконные живут, достигают старости, да и силами крепки?
JOB|21|8|Дети их с ними перед лицем их, и внуки их перед глазами их.
JOB|21|9|Домы их безопасны от страха, и нет жезла Божия на них.
JOB|21|10|Вол их оплодотворяет и не извергает, корова их зачинает и не выкидывает.
JOB|21|11|Как стадо, выпускают они малюток своих, и дети их прыгают.
JOB|21|12|Восклицают под [голос] тимпана и цитры и веселятся при звуках свирели;
JOB|21|13|проводят дни свои в счастьи и мгновенно нисходят в преисподнюю.
JOB|21|14|А между тем они говорят Богу: отойди от нас, не хотим мы знать путей Твоих!
JOB|21|15|Что Вседержитель, чтобы нам служить Ему? и что пользы прибегать к Нему?
JOB|21|16|Видишь, счастье их не от их рук. – Совет нечестивых будь далек от меня!
JOB|21|17|Часто ли угасает светильник у беззаконных, и находит на них беда, и Он дает им в удел страдания во гневе Своем?
JOB|21|18|Они должны быть, как соломинка пред ветром и как плева, уносимая вихрем.
JOB|21|19|[Скажешь]: Бог бережет для детей его несчастье его. – Пусть воздаст Он ему самому, чтобы он это знал.
JOB|21|20|Пусть его глаза увидят несчастье его, и пусть он сам пьет от гнева Вседержителева.
JOB|21|21|Ибо какая ему забота до дома своего после него, когда число месяцев его кончится?
JOB|21|22|Но Бога ли учить мудрости, когда Он судит и горних?
JOB|21|23|Один умирает в самой полноте сил своих, совершенно спокойный и мирный;
JOB|21|24|внутренности его полны жира, и кости его напоены мозгом.
JOB|21|25|А другой умирает с душею огорченною, не вкусив добра.
JOB|21|26|И они вместе будут лежать во прахе, и червь покроет их.
JOB|21|27|Знаю я ваши мысли и ухищрения, какие вы против меня сплетаете.
JOB|21|28|Вы скажете: где дом князя, и где шатер, в котором жили беззаконные?
JOB|21|29|Разве вы не спрашивали у путешественников и незнакомы с их наблюдениями,
JOB|21|30|что в день погибели пощажен бывает злодей, в день гнева отводится в сторону?
JOB|21|31|Кто представит ему пред лице путь его, и кто воздаст ему за то, что он делал?
JOB|21|32|Его провожают ко гробам и на его могиле ставят стражу.
JOB|21|33|Сладки для него глыбы долины, и за ним идет толпа людей, а идущим перед ним нет числа.
JOB|21|34|Как же вы хотите утешать меня пустым? В ваших ответах остается [одна] ложь.
JOB|22|1|И отвечал Елифаз Феманитянин и сказал:
JOB|22|2|разве может человек доставлять пользу Богу? Разумный доставляет пользу себе самому.
JOB|22|3|Что за удовольствие Вседержителю, что ты праведен? И будет ли Ему выгода от того, что ты содержишь пути твои в непорочности?
JOB|22|4|Неужели Он, боясь тебя, вступит с тобою в состязание, пойдет судиться с тобою?
JOB|22|5|Верно, злоба твоя велика, и беззакониям твоим нет конца.
JOB|22|6|Верно, ты брал залоги от братьев твоих ни за что и с полунагих снимал одежду.
JOB|22|7|Утомленному жаждою не подавал воды напиться и голодному отказывал в хлебе;
JOB|22|8|а человеку сильному ты [давал] землю, и сановитый селился на ней.
JOB|22|9|Вдов ты отсылал ни с чем и сирот оставлял с пустыми руками.
JOB|22|10|За то вокруг тебя петли, и возмутил тебя неожиданный ужас,
JOB|22|11|или тьма, в которой ты ничего не видишь, и множество вод покрыло тебя.
JOB|22|12|Не превыше ли небес Бог? посмотри вверх на звезды, как они высоко!
JOB|22|13|И ты говоришь: что знает Бог? может ли Он судить сквозь мрак?
JOB|22|14|Облака – завеса Его, так что Он не видит, а ходит [только] по небесному кругу.
JOB|22|15|Неужели ты держишься пути древних, по которому шли люди беззаконные,
JOB|22|16|которые преждевременно были истреблены, когда вода разлилась под основание их?
JOB|22|17|Они говорили Богу: отойди от нас! и что сделает им Вседержитель?
JOB|22|18|А Он наполнял домы их добром. Но совет нечестивых будь далек от меня!
JOB|22|19|Видели праведники и радовались, и непорочный смеялся им:
JOB|22|20|враг наш истреблен, а оставшееся после них пожрал огонь.
JOB|22|21|Сблизься же с Ним – и будешь спокоен; чрез это придет к тебе добро.
JOB|22|22|Прими из уст Его закон и положи слова Его в сердце твое.
JOB|22|23|Если ты обратишься к Вседержителю, то вновь устроишься, удалишь беззаконие от шатра твоего
JOB|22|24|и будешь вменять в прах блестящий металл, и в камни потоков – [золото] Офирское.
JOB|22|25|И будет Вседержитель твоим золотом и блестящим серебром у тебя,
JOB|22|26|ибо тогда будешь радоваться о Вседержителе и поднимешь к Богу лице твое.
JOB|22|27|Помолишься Ему, и Он услышит тебя, и ты исполнишь обеты твои.
JOB|22|28|Положишь намерение, и оно состоится у тебя, и над путями твоими будет сиять свет.
JOB|22|29|Когда кто уничижен будет, ты скажешь: возвышение! и Он спасет поникшего лицем,
JOB|22|30|избавит и небезвинного, и он спасется чистотою рук твоих.
JOB|23|1|И отвечал Иов и сказал:
JOB|23|2|еще и ныне горька речь моя: страдания мои тяжелее стонов моих.
JOB|23|3|О, если бы я знал, где найти Его, и мог подойти к престолу Его!
JOB|23|4|Я изложил бы пред Ним дело мое и уста мои наполнил бы оправданиями;
JOB|23|5|узнал бы слова, какими Он ответит мне, и понял бы, что Он скажет мне.
JOB|23|6|Неужели Он в полном могуществе стал бы состязаться со мною? О, нет! Пусть Он только обратил бы внимание на меня.
JOB|23|7|Тогда праведник мог бы состязаться с Ним, – и я навсегда получил бы свободу от Судии моего.
JOB|23|8|Но вот, я иду вперед – и нет Его, назад – и не нахожу Его;
JOB|23|9|делает ли Он что на левой стороне, я не вижу; скрывается ли на правой, не усматриваю.
JOB|23|10|Но Он знает путь мой; пусть испытает меня, – выйду, как золото.
JOB|23|11|Нога моя твердо держится стези Его; пути Его я хранил и не уклонялся.
JOB|23|12|От заповеди уст Его не отступал; глаголы уст Его хранил больше, нежели мои правила.
JOB|23|13|Но Он тверд; и кто отклонит Его? Он делает, чего хочет душа Его.
JOB|23|14|Так, Он выполнит положенное мне, и подобного этому много у Него.
JOB|23|15|Поэтому я трепещу пред лицем Его; размышляю – и страшусь Его.
JOB|23|16|Бог расслабил сердце мое, и Вседержитель устрашил меня.
JOB|23|17|Зачем я не уничтожен прежде этой тьмы, и Он не сокрыл мрака от лица моего!
JOB|24|1|Почему не сокрыты от Вседержителя времена, и знающие Его не видят дней Его?
JOB|24|2|Межи передвигают, угоняют стада и пасут [у себя].
JOB|24|3|У сирот уводят осла, у вдовы берут в залог вола;
JOB|24|4|бедных сталкивают с дороги, все уничиженные земли принуждены скрываться.
JOB|24|5|Вот они, [как] дикие ослы в пустыне, выходят на дело свое, вставая рано на добычу; степь [дает] хлеб для них и для детей их;
JOB|24|6|жнут они на поле не своем и собирают виноград у нечестивца;
JOB|24|7|нагие ночуют без покрова и без одеяния на стуже;
JOB|24|8|мокнут от горных дождей и, не имея убежища, жмутся к скале;
JOB|24|9|отторгают от сосцов сироту и с нищего берут залог;
JOB|24|10|заставляют ходить нагими, без одеяния, и голодных кормят колосьями;
JOB|24|11|между стенами выжимают масло оливковое, топчут в точилах и жаждут.
JOB|24|12|В городе люди стонут, и душа убиваемых вопит, и Бог не воспрещает того.
JOB|24|13|Есть из них враги света, не знают путей его и не ходят по стезям его.
JOB|24|14|С рассветом встает убийца, умерщвляет бедного и нищего, а ночью бывает вором.
JOB|24|15|И око прелюбодея ждет сумерков, говоря: ничей глаз не увидит меня, – и закрывает лице.
JOB|24|16|В темноте подкапываются под домы, которые днем они заметили для себя; не знают света.
JOB|24|17|Ибо для них утро – смертная тень, так как они знакомы с ужасами смертной тени.
JOB|24|18|Легок такой на поверхности воды, проклята часть его на земле, и не смотрит он на дорогу садов виноградных.
JOB|24|19|Засуха и жара поглощают снежную воду: так преисподняя – грешников.
JOB|24|20|Пусть забудет его утроба [матери]; пусть лакомится им червь; пусть не остается о нем память; как дерево, пусть сломится беззаконник,
JOB|24|21|который угнетает бездетную, не рождавшую, и вдове не делает добра.
JOB|24|22|Он и сильных увлекает своею силою; он встает и никто не уверен за жизнь свою.
JOB|24|23|А Он дает ему [все] для безопасности, и он [на то] опирается, и очи Его видят пути их.
JOB|24|24|Поднялись высоко, – и вот, нет их; падают и умирают, как и все, и, как верхушки колосьев, срезываются.
JOB|24|25|Если это не так, – кто обличит меня во лжи и в ничто обратит речь мою?
JOB|25|1|И отвечал Вилдад Савхеянин и сказал:
JOB|25|2|держава и страх у Него; Он творит мир на высотах Своих!
JOB|25|3|Есть ли счет воинствам Его? и над кем не восходит свет Его?
JOB|25|4|И как человеку быть правым пред Богом, и как быть чистым рожденному женщиною?
JOB|25|5|Вот даже луна, и та несветла, и звезды нечисты пред очами Его.
JOB|25|6|Тем менее человек, [который] есть червь, и сын человеческий, [который] есть моль.
JOB|26|1|И отвечал Иов и сказал:
JOB|26|2|как ты помог бессильному, поддержал мышцу немощного!
JOB|26|3|Какой совет подал ты немудрому и как во всей полноте объяснил дело!
JOB|26|4|Кому ты говорил эти слова, и чей дух исходил из тебя?
JOB|26|5|Рефаимы трепещут под водами, и живущие в них.
JOB|26|6|Преисподняя обнажена пред Ним, и нет покрывала Аваддону.
JOB|26|7|Он распростер север над пустотою, повесил землю ни на чем.
JOB|26|8|Он заключает воды в облаках Своих, и облако не расседается под ними.
JOB|26|9|Он поставил престол Свой, распростер над ним облако Свое.
JOB|26|10|Черту провел над поверхностью воды, до границ света со тьмою.
JOB|26|11|Столпы небес дрожат и ужасаются от грозы Его.
JOB|26|12|Силою Своею волнует море и разумом Своим сражает его дерзость.
JOB|26|13|От духа Его – великолепие неба; рука Его образовала быстрого скорпиона.
JOB|26|14|Вот, это части путей Его; и как мало мы слышали о Нем! А гром могущества Его кто может уразуметь?
JOB|27|1|И продолжал Иов возвышенную речь свою и сказал:
JOB|27|2|жив Бог, лишивший [меня] суда, и Вседержитель, огорчивший душу мою,
JOB|27|3|что, доколе еще дыхание мое во мне и дух Божий в ноздрях моих,
JOB|27|4|не скажут уста мои неправды, и язык мой не произнесет лжи!
JOB|27|5|Далек я от того, чтобы признать вас справедливыми; доколе не умру, не уступлю непорочности моей.
JOB|27|6|Крепко держал я правду мою и не опущу ее; не укорит меня сердце мое во все дни мои.
JOB|27|7|Враг мой будет, как нечестивец, и восстающий на меня, как беззаконник.
JOB|27|8|Ибо какая надежда лицемеру, когда возьмет, когда исторгнет Бог душу его?
JOB|27|9|Услышит ли Бог вопль его, когда придет на него беда?
JOB|27|10|Будет ли он утешаться Вседержителем и призывать Бога во всякое время?
JOB|27|11|Возвещу вам, что в руке Божией; что у Вседержителя, не скрою.
JOB|27|12|Вот, все вы и сами видели; и для чего вы столько пустословите?
JOB|27|13|Вот доля человеку беззаконному от Бога, и наследие, какое получают от Вседержителя притеснители.
JOB|27|14|Если умножаются сыновья его, то под меч; и потомки его не насытятся хлебом.
JOB|27|15|Оставшихся по нем смерть низведет во гроб, и вдовы их не будут плакать.
JOB|27|16|Если он наберет кучи серебра, как праха, и наготовит одежд, как брение,
JOB|27|17|то он наготовит, а одеваться будет праведник, и серебро получит себе на долю беспорочный.
JOB|27|18|Он строит, как моль, дом свой и, как сторож, делает себе шалаш;
JOB|27|19|ложится спать богачом и таким не встанет; открывает глаза свои, и он уже не тот.
JOB|27|20|Как воды, постигнут его ужасы; в ночи похитит его буря.
JOB|27|21|Поднимет его восточный ветер и понесет, и он быстро побежит от него.
JOB|27|22|Устремится на него и не пощадит, как бы он ни силился убежать от руки его.
JOB|27|23|Всплеснут о нем руками и посвищут над ним с места его!
JOB|28|1|Так! у серебра есть источная жила, и у золота место, [где его] плавят.
JOB|28|2|Железо получается из земли; из камня выплавляется медь.
JOB|28|3|[Человек] полагает предел тьме и тщательно разыскивает камень во мраке и тени смертной.
JOB|28|4|Вырывают рудокопный колодезь в местах, забытых ногою, спускаются вглубь, висят [и] зыблются вдали от людей.
JOB|28|5|Земля, на которой вырастает хлеб, внутри изрыта как бы огнем.
JOB|28|6|Камни ее – место сапфира, и в ней песчинки золота.
JOB|28|7|Стези [туда] не знает хищная птица, и не видал ее глаз коршуна;
JOB|28|8|не попирали ее скимны, и не ходил по ней шакал.
JOB|28|9|На гранит налагает он руку свою, с корнем опрокидывает горы;
JOB|28|10|в скалах просекает каналы, и все драгоценное видит глаз его;
JOB|28|11|останавливает течение потоков и сокровенное выносит на свет.
JOB|28|12|Но где премудрость обретается? и где место разума?
JOB|28|13|Не знает человек цены ее, и она не обретается на земле живых.
JOB|28|14|Бездна говорит: не во мне она; и море говорит: не у меня.
JOB|28|15|Не дается она за золото и не приобретается она за вес серебра;
JOB|28|16|не оценивается она золотом Офирским, ни драгоценным ониксом, ни сапфиром;
JOB|28|17|не равняется с нею золото и кристалл, и не выменяешь ее на сосуды из чистого золота.
JOB|28|18|А о кораллах и жемчуге и упоминать нечего, и приобретение премудрости выше рубинов.
JOB|28|19|Не равняется с нею топаз Ефиопский; чистым золотом не оценивается она.
JOB|28|20|Откуда же исходит премудрость? и где место разума?
JOB|28|21|Сокрыта она от очей всего живущего и от птиц небесных утаена.
JOB|28|22|Аваддон и смерть говорят: ушами нашими слышали мы слух о ней.
JOB|28|23|Бог знает путь ее, и Он ведает место ее.
JOB|28|24|Ибо Он прозирает до концов земли и видит под всем небом.
JOB|28|25|Когда Он ветру полагал вес и располагал воду по мере,
JOB|28|26|когда назначал устав дождю и путь для молнии громоносной,
JOB|28|27|тогда Он видел ее и явил ее, приготовил ее и еще испытал ее
JOB|28|28|и сказал человеку: вот, страх Господень есть истинная премудрость, и удаление от зла – разум.
JOB|29|1|И продолжал Иов возвышенную речь свою и сказал:
JOB|29|2|о, если бы я был, как в прежние месяцы, как в те дни, когда Бог хранил меня,
JOB|29|3|когда светильник Его светил над головою моею, и я при свете Его ходил среди тьмы;
JOB|29|4|как был я во дни молодости моей, когда милость Божия [была] над шатром моим,
JOB|29|5|когда еще Вседержитель [был] со мною, и дети мои вокруг меня,
JOB|29|6|когда пути мои обливались молоком, и скала источала для меня ручьи елея!
JOB|29|7|когда я выходил к воротам города и на площади ставил седалище свое, –
JOB|29|8|юноши, увидев меня, прятались, а старцы вставали и стояли;
JOB|29|9|князья удерживались от речи и персты полагали на уста свои;
JOB|29|10|голос знатных умолкал, и язык их прилипал к гортани их.
JOB|29|11|Ухо, слышавшее меня, ублажало меня; око видевшее восхваляло меня,
JOB|29|12|потому что я спасал страдальца вопиющего и сироту беспомощного.
JOB|29|13|Благословение погибавшего приходило на меня, и сердцу вдовы доставлял я радость.
JOB|29|14|Я облекался в правду, и суд мой одевал меня, как мантия и увясло.
JOB|29|15|Я был глазами слепому и ногами хромому;
JOB|29|16|отцом был я для нищих и тяжбу, которой я не знал, разбирал внимательно.
JOB|29|17|Сокрушал я беззаконному челюсти и из зубов его исторгал похищенное.
JOB|29|18|И говорил я: в гнезде моем скончаюсь, и дни [мои] будут многи, как песок;
JOB|29|19|корень мой открыт для воды, и роса ночует на ветвях моих;
JOB|29|20|слава моя не стареет, лук мой крепок в руке моей.
JOB|29|21|Внимали мне и ожидали, и безмолвствовали при совете моем.
JOB|29|22|После слов моих уже не рассуждали; речь моя капала на них.
JOB|29|23|Ждали меня, как дождя, и, [как] дождю позднему, открывали уста свои.
JOB|29|24|Бывало, улыбнусь им – они не верят; и света лица моего они не помрачали.
JOB|29|25|Я назначал пути им и сидел во главе и жил как царь в кругу воинов, как утешитель плачущих.
JOB|30|1|А ныне смеются надо мною младшие меня летами, те, которых отцов я не согласился бы поместить с псами стад моих.
JOB|30|2|И сила рук их к чему мне? Над ними уже прошло время.
JOB|30|3|Бедностью и голодом истощенные, они убегают в степь безводную, мрачную и опустевшую;
JOB|30|4|щиплют зелень подле кустов, и ягоды можжевельника – хлеб их.
JOB|30|5|Из общества изгоняют их, кричат на них, как на воров,
JOB|30|6|чтобы жили они в рытвинах потоков, в ущельях земли и утесов.
JOB|30|7|Ревут между кустами, жмутся под терном.
JOB|30|8|Люди отверженные, люди без имени, отребье земли!
JOB|30|9|Их–то сделался я ныне песнью и пищею разговора их.
JOB|30|10|Они гнушаются мною, удаляются от меня и не удерживаются плевать пред лицем моим.
JOB|30|11|Так как Он развязал повод мой и поразил меня, то они сбросили с себя узду пред лицем моим.
JOB|30|12|С правого боку встает это исчадие, сбивает меня с ног, направляет гибельные свои пути ко мне.
JOB|30|13|А мою стезю испортили: все успели сделать к моей погибели, не имея помощника.
JOB|30|14|Они пришли ко мне, как сквозь широкий пролом; с шумом бросились на меня.
JOB|30|15|Ужасы устремились на меня; как ветер, развеялось величие мое, и счастье мое унеслось, как облако.
JOB|30|16|И ныне изливается душа моя во мне: дни скорби объяли меня.
JOB|30|17|Ночью ноют во мне кости мои, и жилы мои не имеют покоя.
JOB|30|18|С великим трудом снимается с меня одежда моя; края хитона моего жмут меня.
JOB|30|19|Он бросил меня в грязь, и я стал, как прах и пепел.
JOB|30|20|Я взываю к Тебе, и Ты не внимаешь мне, – стою, а Ты [только] смотришь на меня.
JOB|30|21|Ты сделался жестоким ко мне, крепкою рукою враждуешь против меня.
JOB|30|22|Ты поднял меня и заставил меня носиться по ветру и сокрушаешь меня.
JOB|30|23|Так, я знаю, что Ты приведешь меня к смерти и в дом собрания всех живущих.
JOB|30|24|Верно, Он не прострет руки Своей на дом костей: будут ли они кричать при своем разрушении?
JOB|30|25|Не плакал ли я о том, кто был в горе? не скорбела ли душа моя о бедных?
JOB|30|26|Когда я чаял добра, пришло зло; когда ожидал света, пришла тьма.
JOB|30|27|Мои внутренности кипят и не перестают; встретили меня дни печали.
JOB|30|28|Я хожу почернелый, но не от солнца; встаю в собрании и кричу.
JOB|30|29|Я стал братом шакалам и другом страусам.
JOB|30|30|Моя кожа почернела на мне, и кости мои обгорели от жара.
JOB|30|31|И цитра моя сделалась унылою, и свирель моя – голосом плачевным.
JOB|31|1|Завет положил я с глазами моими, чтобы не помышлять мне о девице.
JOB|31|2|Какая же участь [мне] от Бога свыше? И какое наследие от Вседержителя с небес?
JOB|31|3|Не для нечестивого ли гибель, и не для делающего ли зло напасть?
JOB|31|4|Не видел ли Он путей моих, и не считал ли всех моих шагов?
JOB|31|5|Если я ходил в суете, и если нога моя спешила на лукавство, –
JOB|31|6|пусть взвесят меня на весах правды, и Бог узнает мою непорочность.
JOB|31|7|Если стопы мои уклонялись от пути и сердце мое следовало за глазами моими, и если что–либо нечистое пристало к рукам моим,
JOB|31|8|то пусть я сею, а другой ест, и пусть отрасли мои искоренены будут.
JOB|31|9|Если сердце мое прельщалось женщиною и я строил ковы у дверей моего ближнего, –
JOB|31|10|пусть моя жена мелет на другого, и пусть другие издеваются над нею,
JOB|31|11|потому что это – преступление, это – беззаконие, подлежащее суду;
JOB|31|12|это – огонь, поядающий до истребления, который искоренил бы все добро мое.
JOB|31|13|Если я пренебрегал правами слуги и служанки моей, когда они имели спор со мною,
JOB|31|14|то что стал бы я делать, когда бы Бог восстал? И когда бы Он взглянул на меня, что мог бы я отвечать Ему?
JOB|31|15|Не Он ли, Который создал меня во чреве, создал и его и равно образовал нас в утробе?
JOB|31|16|Отказывал ли я нуждающимся в их просьбе и томил ли глаза вдовы?
JOB|31|17|Один ли я съедал кусок мой, и не ел ли от него и сирота?
JOB|31|18|Ибо с детства он рос со мною, как с отцом, и от чрева матери моей я руководил [вдову].
JOB|31|19|Если я видел кого погибавшим без одежды и бедного без покрова, –
JOB|31|20|не благословляли ли меня чресла его, и не был ли он согрет шерстью овец моих?
JOB|31|21|Если я поднимал руку мою на сироту, когда видел помощь себе у ворот,
JOB|31|22|то пусть плечо мое отпадет от спины, и рука моя пусть отломится от локтя,
JOB|31|23|ибо страшно для меня наказание от Бога: пред величием Его не устоял бы я.
JOB|31|24|Полагал ли я в золоте опору мою и говорил ли сокровищу: ты – надежда моя?
JOB|31|25|Радовался ли я, что богатство мое было велико, и что рука моя приобрела много?
JOB|31|26|Смотря на солнце, как оно сияет, и на луну, как она величественно шествует,
JOB|31|27|прельстился ли я в тайне сердца моего, и целовали ли уста мои руку мою?
JOB|31|28|Это также было бы преступление, подлежащее суду, потому что я отрекся бы [тогда] от Бога Всевышнего.
JOB|31|29|Радовался ли я погибели врага моего и торжествовал ли, когда несчастье постигало его?
JOB|31|30|Не позволял я устам моим грешить проклятием души его.
JOB|31|31|Не говорили ли люди шатра моего: о, если бы мы от мяс его не насытились?
JOB|31|32|Странник не ночевал на улице; двери мои я отворял прохожему.
JOB|31|33|Если бы я скрывал проступки мои, как человек, утаивая в груди моей пороки мои,
JOB|31|34|то я боялся бы большого общества, и презрение одноплеменников страшило бы меня, и я молчал бы и не выходил бы за двери.
JOB|31|35|О, если бы кто выслушал меня! Вот мое желание, чтобы Вседержитель отвечал мне, и чтобы защитник мой составил запись.
JOB|31|36|Я носил бы ее на плечах моих и возлагал бы ее, как венец;
JOB|31|37|объявил бы ему число шагов моих, сблизился бы с ним, как с князем.
JOB|31|38|Если вопияла на меня земля моя и жаловались на меня борозды ее;
JOB|31|39|если я ел плоды ее без платы и отягощал жизнь земледельцев,
JOB|31|40|то пусть вместо пшеницы вырастает волчец и вместо ячменя куколь. Слова Иова кончились.
JOB|32|1|Когда те три мужа перестали отвечать Иову, потому что он был прав в глазах своих,
JOB|32|2|тогда воспылал гнев Елиуя, сына Варахиилова, Вузитянина из племени Рамова: воспылал гнев его на Иова за то, что он оправдывал себя больше, нежели Бога,
JOB|32|3|а на трех друзей его воспылал гнев его за то, что они не нашли, что отвечать, а между тем обвиняли Иова.
JOB|32|4|Елиуй ждал, пока Иов говорил, потому что они летами были старше его.
JOB|32|5|Когда же Елиуй увидел, что нет ответа в устах тех трех мужей, тогда воспылал гнев его.
JOB|32|6|И отвечал Елиуй, сын Варахиилов, Вузитянин, и сказал: я молод летами, а вы – старцы; поэтому я робел и боялся объявлять вам мое мнение.
JOB|32|7|Я говорил сам себе: пусть говорят дни, и многолетие поучает мудрости.
JOB|32|8|Но дух в человеке и дыхание Вседержителя дает ему разумение.
JOB|32|9|Не многолетние [только] мудры, и не старики разумеют правду.
JOB|32|10|Поэтому я говорю: выслушайте меня, объявлю вам мое мнение и я.
JOB|32|11|Вот, я ожидал слов ваших, – вслушивался в суждения ваши, доколе вы придумывали, что сказать.
JOB|32|12|Я пристально смотрел на вас, и вот никто из вас не обличает Иова и не отвечает на слова его.
JOB|32|13|Не скажите: мы нашли мудрость: Бог опровергнет его, а не человек.
JOB|32|14|Если бы он обращал слова свои ко мне, то я не вашими речами отвечал бы ему.
JOB|32|15|Испугались, не отвечают более; перестали говорить.
JOB|32|16|И как я ждал, а они не говорят, остановились и не отвечают более,
JOB|32|17|то и я отвечу с моей стороны, объявлю мое мнение и я,
JOB|32|18|ибо я полон речами, и дух во мне теснит меня.
JOB|32|19|Вот, утроба моя, как вино неоткрытое: она готова прорваться, подобно новым мехам.
JOB|32|20|Поговорю, и будет легче мне; открою уста мои и отвечу.
JOB|32|21|На лице человека смотреть не буду и никакому человеку льстить не стану,
JOB|32|22|потому что я не умею льстить: сейчас убей меня, Творец мой.
JOB|33|1|Итак слушай, Иов, речи мои и внимай всем словам моим.
JOB|33|2|Вот, я открываю уста мои, язык мой говорит в гортани моей.
JOB|33|3|Слова мои от искренности моего сердца, и уста мои произнесут знание чистое.
JOB|33|4|Дух Божий создал меня, и дыхание Вседержителя дало мне жизнь.
JOB|33|5|Если можешь, отвечай мне и стань передо мною.
JOB|33|6|Вот я, по желанию твоему, вместо Бога. Я образован также из брения;
JOB|33|7|поэтому страх передо мною не может смутить тебя, и рука моя не будет тяжела для тебя.
JOB|33|8|Ты говорил в уши мои, и я слышал звук слов:
JOB|33|9|чист я, без порока, невинен я, и нет во мне неправды;
JOB|33|10|а Он нашел обвинение против меня и считает меня Своим противником;
JOB|33|11|поставил ноги мои в колоду, наблюдает за всеми путями моими.
JOB|33|12|Вот в этом ты неправ, отвечаю тебе, потому что Бог выше человека.
JOB|33|13|Для чего тебе состязаться с Ним? Он не дает отчета ни в каких делах Своих.
JOB|33|14|Бог говорит однажды и, если того не заметят, в другой раз:
JOB|33|15|во сне, в ночном видении, когда сон находит на людей, во время дремоты на ложе.
JOB|33|16|Тогда Он открывает у человека ухо и запечатлевает Свое наставление,
JOB|33|17|чтобы отвести человека от какого–либо предприятия и удалить от него гордость,
JOB|33|18|чтобы отвести душу его от пропасти и жизнь его от поражения мечом.
JOB|33|19|Или он вразумляется болезнью на ложе своем и жестокою болью во всех костях своих, –
JOB|33|20|и жизнь его отвращается от хлеба и душа его от любимой пищи.
JOB|33|21|Плоть на нем пропадает, так что ее не видно, и показываются кости его, которых не было видно.
JOB|33|22|И душа его приближается к могиле и жизнь его – к смерти.
JOB|33|23|Если есть у него Ангел–наставник, один из тысячи, чтобы показать человеку прямой [путь] его, –
JOB|33|24|[Бог] умилосердится над ним и скажет: освободи его от могилы; Я нашел умилостивление.
JOB|33|25|Тогда тело его сделается свежее, нежели в молодости; он возвратится к дням юности своей.
JOB|33|26|Будет молиться Богу, и Он – милостив к нему; с радостью взирает на лице его и возвращает человеку праведность его.
JOB|33|27|Он будет смотреть на людей и говорить: грешил я и превращал правду, и не воздано мне;
JOB|33|28|Он освободил душу мою от могилы, и жизнь моя видит свет.
JOB|33|29|Вот, все это делает Бог два–три раза с человеком,
JOB|33|30|чтобы отвести душу его от могилы и просветить его светом живых.
JOB|33|31|Внимай, Иов, слушай меня, молчи, и я буду говорить.
JOB|33|32|Если имеешь, что сказать, отвечай; говори, потому что я желал бы твоего оправдания;
JOB|33|33|если же нет, то слушай меня: молчи, и я научу тебя мудрости.
JOB|34|1|И продолжал Елиуй и сказал:
JOB|34|2|выслушайте, мудрые, речь мою, и приклоните ко мне ухо, рассудительные!
JOB|34|3|Ибо ухо разбирает слова, как гортань различает вкус в пище.
JOB|34|4|Установим между собою рассуждение и распознаем, что хорошо.
JOB|34|5|Вот, Иов сказал: я прав, но Бог лишил меня суда.
JOB|34|6|Должен ли я лгать на правду мою? Моя рана неисцелима без вины.
JOB|34|7|Есть ли такой человек, как Иов, который пьет глумление, как воду,
JOB|34|8|вступает в сообщество с делающими беззаконие и ходит с людьми нечестивыми?
JOB|34|9|Потому что он сказал: нет пользы для человека в благоугождении Богу.
JOB|34|10|Итак послушайте меня, мужи мудрые! Не может быть у Бога неправда или у Вседержителя неправосудие,
JOB|34|11|ибо Он по делам человека поступает с ним и по путям мужа воздает ему.
JOB|34|12|Истинно, Бог не делает неправды и Вседержитель не извращает суда.
JOB|34|13|Кто кроме Его промышляет о земле? И кто управляет всею вселенною?
JOB|34|14|Если бы Он обратил сердце Свое к Себе и взял к Себе дух ее и дыхание ее, –
JOB|34|15|вдруг погибла бы всякая плоть, и человек возвратился бы в прах.
JOB|34|16|Итак, если ты имеешь разум, то слушай это и внимай словам моим.
JOB|34|17|Ненавидящий правду может ли владычествовать? И можешь ли ты обвинить Всеправедного?
JOB|34|18|Можно ли сказать царю: ты – нечестивец, и князьям: вы – беззаконники?
JOB|34|19|Но Он не смотрит и на лица князей и не предпочитает богатого бедному, потому что все они дело рук Его.
JOB|34|20|Внезапно они умирают; среди ночи народ возмутится, и они исчезают; и сильных изгоняют не силою.
JOB|34|21|Ибо очи Его над путями человека, и Он видит все шаги его.
JOB|34|22|Нет тьмы, ни тени смертной, где могли бы укрыться делающие беззаконие.
JOB|34|23|Потому Он уже не требует от человека, чтобы шел на суд с Богом.
JOB|34|24|Он сокрушает сильных без исследования и поставляет других на их места;
JOB|34|25|потому что Он делает известными дела их и низлагает их ночью, и они истребляются.
JOB|34|26|Он поражает их, как беззаконных людей, пред глазами других,
JOB|34|27|за то, что они отвратились от Него и не уразумели всех путей Его,
JOB|34|28|так что дошел до Него вопль бедных, и Он услышал стенание угнетенных.
JOB|34|29|Дарует ли Он тишину, кто может возмутить? скрывает ли Он лице Свое, кто может увидеть Его? Будет ли это для народа, или для одного человека,
JOB|34|30|чтобы не царствовал лицемер к соблазну народа.
JOB|34|31|К Богу должно говорить: я потерпел, больше не буду грешить.
JOB|34|32|А чего я не знаю, Ты научи меня; и если я сделал беззаконие, больше не буду.
JOB|34|33|По твоему ли [рассуждению] Он должен воздавать? И как ты отвергаешь, то тебе следует избирать, а не мне; говори, что знаешь.
JOB|34|34|Люди разумные скажут мне, и муж мудрый, слушающий меня:
JOB|34|35|Иов не умно говорит, и слова его не со смыслом.
JOB|34|36|Я желал бы, чтобы Иов вполне был испытан, по ответам его, свойственным людям нечестивым.
JOB|34|37|Иначе он ко греху своему прибавит отступление, будет рукоплескать между нами и еще больше наговорит против Бога.
JOB|35|1|И продолжал Елиуй и сказал:
JOB|35|2|считаешь ли ты справедливым, что сказал: я правее Бога?
JOB|35|3|Ты сказал: что пользы мне? и какую прибыль я имел бы пред тем, как если бы я и грешил?
JOB|35|4|Я отвечу тебе и твоим друзьям с тобою:
JOB|35|5|взгляни на небо и смотри; воззри на облака, они выше тебя.
JOB|35|6|Если ты грешишь, что делаешь ты Ему? и если преступления твои умножаются, что причиняешь ты Ему?
JOB|35|7|Если ты праведен, что даешь Ему? или что получает Он от руки твоей?
JOB|35|8|Нечестие твое относится к человеку, как ты, и праведность твоя к сыну человеческому.
JOB|35|9|От множества притеснителей стонут притесняемые, и от руки сильных вопиют.
JOB|35|10|Но никто не говорит: где Бог, Творец мой, Который дает песни в ночи,
JOB|35|11|Который научает нас более, нежели скотов земных, и вразумляет нас более, нежели птиц небесных?
JOB|35|12|Там они вопиют, и Он не отвечает им, по причине гордости злых людей.
JOB|35|13|Но неправда, что Бог не слышит и Вседержитель не взирает на это.
JOB|35|14|Хотя ты сказал, что ты не видишь Его, но суд пред Ним, и – жди его.
JOB|35|15|Но ныне, потому что гнев Его не посетил его и он не познал его во всей строгости,
JOB|35|16|Иов и открыл легкомысленно уста свои и безрассудно расточает слова.
JOB|36|1|И продолжал Елиуй и сказал:
JOB|36|2|подожди меня немного, и я покажу тебе, что я имею еще что сказать за Бога.
JOB|36|3|Начну мои рассуждения издалека и воздам Создателю моему справедливость,
JOB|36|4|потому что слова мои точно не ложь: пред тобою – совершенный в познаниях.
JOB|36|5|Вот, Бог могуществен и не презирает сильного крепостью сердца;
JOB|36|6|Он не поддерживает нечестивых и воздает должное угнетенным;
JOB|36|7|Он не отвращает очей Своих от праведников, но с царями навсегда посаждает их на престоле, и они возвышаются.
JOB|36|8|Если же они окованы цепями и содержатся в узах бедствия,
JOB|36|9|то Он указывает им на дела их и на беззакония их, потому что умножились,
JOB|36|10|и открывает их ухо для вразумления и говорит им, чтоб они отстали от нечестия.
JOB|36|11|Если послушают и будут служить Ему, то проведут дни свои в благополучии и лета свои в радости;
JOB|36|12|если же не послушают, то погибнут от стрелы и умрут в неразумии.
JOB|36|13|Но лицемеры питают в сердце гнев и не взывают к Нему, когда Он заключает их в узы;
JOB|36|14|поэтому душа их умирает в молодости и жизнь их с блудниками.
JOB|36|15|Он спасает бедного от беды его и в угнетении открывает ухо его.
JOB|36|16|И тебя вывел бы Он из тесноты на простор, где нет стеснения, и поставляемое на стол твой было бы наполнено туком;
JOB|36|17|но ты преисполнен суждениями нечестивых: суждение и осуждение – близки.
JOB|36|18|Да не поразит тебя гнев [Божий] наказанием! Большой выкуп не спасет тебя.
JOB|36|19|Даст ли Он какую цену твоему богатству? Нет, – ни золоту и никакому сокровищу.
JOB|36|20|Не желай той ночи, когда народы истребляются на своем месте.
JOB|36|21|Берегись, не склоняйся к нечестию, которое ты предпочел страданию.
JOB|36|22|Бог высок могуществом Своим, и кто такой, как Он, наставник?
JOB|36|23|Кто укажет Ему путь Его; кто может сказать: Ты поступаешь несправедливо?
JOB|36|24|Помни о том, чтобы превозносить дела его, которые люди видят.
JOB|36|25|Все люди могут видеть их; человек может усматривать их издали.
JOB|36|26|Вот, Бог велик, и мы не можем познать Его; число лет Его неисследимо.
JOB|36|27|Он собирает капли воды; они во множестве изливаются дождем:
JOB|36|28|из облаков каплют и изливаются обильно на людей.
JOB|36|29|Кто может также постигнуть протяжение облаков, треск шатра Его?
JOB|36|30|Вот, Он распространяет над ним свет Свой и покрывает дно моря.
JOB|36|31|Оттуда Он судит народы, дает пищу в изобилии.
JOB|36|32|Он сокрывает в дланях Своих молнию и повелевает ей, кого разить.
JOB|36|33|Треск ее дает знать о ней; скот также чувствует происходящее.
JOB|37|1|И от сего трепещет сердце мое и подвиглось с места своего.
JOB|37|2|Слушайте, слушайте голос Его и гром, исходящий из уст Его.
JOB|37|3|Под всем небом раскат его, и блистание его – до краев земли.
JOB|37|4|За ним гремит глас; гремит Он гласом величества Своего и не останавливает его, когда голос Его услышан.
JOB|37|5|Дивно гремит Бог гласом Своим, делает дела великие, для нас непостижимые.
JOB|37|6|Ибо снегу Он говорит: будь на земле; равно мелкий дождь и большой дождь в Его власти.
JOB|37|7|Он полагает печать на руку каждого человека, чтобы все люди знали дело Его.
JOB|37|8|Тогда зверь уходит в убежище и остается в своих логовищах.
JOB|37|9|От юга приходит буря, от севера – стужа.
JOB|37|10|От дуновения Божия происходит лед, и поверхность воды сжимается.
JOB|37|11|Также влагою Он наполняет тучи, и облака сыплют свет Его,
JOB|37|12|и они направляются по намерениям Его, чтоб исполнить то, что Он повелит им на лице обитаемой земли.
JOB|37|13|Он повелевает им идти или для наказания, или в благоволение, или для помилования.
JOB|37|14|Внимай сему, Иов; стой и разумевай чудные дела Божии.
JOB|37|15|Знаешь ли, как Бог располагает ими и повелевает свету блистать из облака Своего?
JOB|37|16|Разумеешь ли равновесие облаков, чудное дело Совершеннейшего в знании?
JOB|37|17|Как нагревается твоя одежда, когда Он успокаивает землю от юга?
JOB|37|18|Ты ли с Ним распростер небеса, твердые, как литое зеркало?
JOB|37|19|Научи нас, что сказать Ему? Мы в этой тьме ничего не можем сообразить.
JOB|37|20|Будет ли возвещено Ему, что я говорю? Сказал ли кто, что сказанное доносится Ему?
JOB|37|21|Теперь не видно яркого света в облаках, но пронесется ветер и расчистит их.
JOB|37|22|Светлая погода приходит от севера, и окрест Бога страшное великолепие.
JOB|37|23|Вседержитель! мы не постигаем Его. Он велик силою, судом и полнотою правосудия. Он [никого] не угнетает.
JOB|37|24|Посему да благоговеют пред Ним люди, и да трепещут пред Ним все мудрые сердцем!
JOB|38|1|Господь отвечал Иову из бури и сказал:
JOB|38|2|кто сей, омрачающий Провидение словами без смысла?
JOB|38|3|Препояшь ныне чресла твои, как муж: Я буду спрашивать тебя, и ты объясняй Мне:
JOB|38|4|где был ты, когда Я полагал основания земли? Скажи, если знаешь.
JOB|38|5|Кто положил меру ей, если знаешь? или кто протягивал по ней вервь?
JOB|38|6|На чем утверждены основания ее, или кто положил краеугольный камень ее,
JOB|38|7|при общем ликовании утренних звезд, когда все сыны Божии восклицали от радости?
JOB|38|8|Кто затворил море воротами, когда оно исторглось, вышло как бы из чрева,
JOB|38|9|когда Я облака сделал одеждою его и мглу пеленами его,
JOB|38|10|и утвердил ему Мое определение, и поставил запоры и ворота,
JOB|38|11|и сказал: доселе дойдешь и не перейдешь, и здесь предел надменным волнам твоим?
JOB|38|12|Давал ли ты когда в жизни своей приказания утру и указывал ли заре место ее,
JOB|38|13|чтобы она охватила края земли и стряхнула с нее нечестивых,
JOB|38|14|чтобы [земля] изменилась, как глина под печатью, и стала, как разноцветная одежда,
JOB|38|15|и чтобы отнялся у нечестивых свет их и дерзкая рука их сокрушилась?
JOB|38|16|Нисходил ли ты во глубину моря и входил ли в исследование бездны?
JOB|38|17|Отворялись ли для тебя врата смерти, и видел ли ты врата тени смертной?
JOB|38|18|Обозрел ли ты широту земли? Объясни, если знаешь все это.
JOB|38|19|Где путь к жилищу света, и где место тьмы?
JOB|38|20|Ты, конечно, доходил до границ ее и знаешь стези к дому ее.
JOB|38|21|Ты знаешь это, потому что ты был уже тогда рожден, и число дней твоих очень велико.
JOB|38|22|Входил ли ты в хранилища снега и видел ли сокровищницы града,
JOB|38|23|которые берегу Я на время смутное, на день битвы и войны?
JOB|38|24|По какому пути разливается свет и разносится восточный ветер по земле?
JOB|38|25|Кто проводит протоки для излияния воды и путь для громоносной молнии,
JOB|38|26|чтобы шел дождь на землю безлюдную, на пустыню, где нет человека,
JOB|38|27|чтобы насыщать пустыню и степь и возбуждать травные зародыши к возрастанию?
JOB|38|28|Есть ли у дождя отец? или кто рождает капли росы?
JOB|38|29|Из чьего чрева выходит лед, и иней небесный, – кто рождает его?
JOB|38|30|Воды, как камень, крепнут, и поверхность бездны замерзает.
JOB|38|31|Можешь ли ты связать узел Хима и разрешить узы Кесиль?
JOB|38|32|Можешь ли выводить созвездия в свое время и вести Ас с ее детьми?
JOB|38|33|Знаешь ли ты уставы неба, можешь ли установить господство его на земле?
JOB|38|34|Можешь ли возвысить голос твой к облакам, чтобы вода в обилии покрыла тебя?
JOB|38|35|Можешь ли посылать молнии, и пойдут ли они и скажут ли тебе: вот мы?
JOB|38|36|Кто вложил мудрость в сердце, или кто дал смысл разуму?
JOB|38|37|Кто может расчислить облака своею мудростью и удержать сосуды неба,
JOB|38|38|когда пыль обращается в грязь и глыбы слипаются?
JOB|38|39|Ты ли ловишь добычу львице и насыщаешь молодых львов,
JOB|38|40|когда они лежат в берлогах или покоятся под тенью в засаде?
JOB|38|41|Кто приготовляет ворону корм его, когда птенцы его кричат к Богу, бродя без пищи?
JOB|39|1|Знаешь ли ты время, когда рождаются дикие козы на скалах, и замечал ли роды ланей?
JOB|39|2|можешь ли расчислить месяцы беременности их? и знаешь ли время родов их?
JOB|39|3|Они изгибаются, рождая детей своих, выбрасывая свои ноши;
JOB|39|4|дети их приходят в силу, растут на поле, уходят и не возвращаются к ним.
JOB|39|5|Кто пустил дикого осла на свободу, и кто разрешил узы онагру,
JOB|39|6|которому степь Я назначил домом и солончаки – жилищем?
JOB|39|7|Он посмевается городскому многолюдству и не слышит криков погонщика,
JOB|39|8|по горам ищет себе пищи и гоняется за всякою зеленью.
JOB|39|9|Захочет ли единорог служить тебе и переночует ли у яслей твоих?
JOB|39|10|Можешь ли веревкою привязать единорога к борозде, и станет ли он боронить за тобою поле?
JOB|39|11|Понадеешься ли на него, потому что у него сила велика, и предоставишь ли ему работу твою?
JOB|39|12|Поверишь ли ему, что он семена твои возвратит и сложит на гумно твое?
JOB|39|13|Ты ли дал красивые крылья павлину и перья и пух страусу?
JOB|39|14|Он оставляет яйца свои на земле, и на песке согревает их,
JOB|39|15|и забывает, что нога может раздавить их и полевой зверь может растоптать их;
JOB|39|16|он жесток к детям своим, как бы не своим, и не опасается, что труд его будет напрасен;
JOB|39|17|потому что Бог не дал ему мудрости и не уделил ему смысла;
JOB|39|18|а когда поднимется на высоту, посмевается коню и всаднику его.
JOB|39|19|Ты ли дал коню силу и облек шею его гривою?
JOB|39|20|Можешь ли ты испугать его, как саранчу? Храпение ноздрей его – ужас;
JOB|39|21|роет ногою землю и восхищается силою; идет навстречу оружию;
JOB|39|22|он смеется над опасностью и не робеет и не отворачивается от меча;
JOB|39|23|колчан звучит над ним, сверкает копье и дротик;
JOB|39|24|в порыве и ярости он глотает землю и не может стоять при звуке трубы;
JOB|39|25|при трубном звуке он издает голос: гу! гу! и издалека чует битву, громкие голоса вождей и крик.
JOB|39|26|Твоею ли мудростью летает ястреб и направляет крылья свои на полдень?
JOB|39|27|По твоему ли слову возносится орел и устрояет на высоте гнездо свое?
JOB|39|28|Он живет на скале и ночует на зубце утесов и на местах неприступных;
JOB|39|29|оттуда высматривает себе пищу: глаза его смотрят далеко;
JOB|39|30|птенцы его пьют кровь, и где труп, там и он.
JOB|40|1|И продолжал Господь и сказал Иову:
JOB|40|2|будет ли состязающийся со Вседержителем еще учить? Обличающий Бога пусть отвечает Ему.
JOB|40|3|И отвечал Иов Господу и сказал:
JOB|40|4|вот, я ничтожен; что буду я отвечать Тебе? Руку мою полагаю на уста мои.
JOB|40|5|Однажды я говорил, – теперь отвечать не буду, даже дважды, но более не буду.
JOB|40|6|И отвечал Господь Иову из бури и сказал:
JOB|40|7|препояшь, как муж, чресла твои: Я буду спрашивать тебя, а ты объясняй Мне.
JOB|40|8|Ты хочешь ниспровергнуть суд Мой, обвинить Меня, чтобы оправдать себя?
JOB|40|9|Такая ли у тебя мышца, как у Бога? И можешь ли возгреметь голосом, как Он?
JOB|40|10|Укрась же себя величием и славою, облекись в блеск и великолепие;
JOB|40|11|излей ярость гнева твоего, посмотри на все гордое и смири его;
JOB|40|12|взгляни на всех высокомерных и унизь их, и сокруши нечестивых на местах их;
JOB|40|13|зарой всех их в землю и лица их покрой тьмою.
JOB|40|14|Тогда и Я признаю, что десница твоя может спасать тебя.
JOB|40|15|Вот бегемот, которого Я создал, как и тебя; он ест траву, как вол;
JOB|40|16|вот, его сила в чреслах его и крепость его в мускулах чрева его;
JOB|40|17|поворачивает хвостом своим, как кедром; жилы же на бедрах его переплетены;
JOB|40|18|ноги у него, как медные трубы; кости у него, как железные прутья;
JOB|40|19|это – верх путей Божиих; только Сотворивший его может приблизить к нему меч Свой;
JOB|40|20|горы приносят ему пищу, и там все звери полевые играют;
JOB|40|21|он ложится под тенистыми деревьями, под кровом тростника и в болотах;
JOB|40|22|тенистые дерева покрывают его своею тенью; ивы при ручьях окружают его;
JOB|40|23|вот, он пьет из реки и не торопится; остается спокоен, хотя бы Иордан устремился ко рту его.
JOB|40|24|Возьмет ли кто его в глазах его и проколет ли ему нос багром?
JOB|40|25|Можешь ли ты удою вытащить левиафана и веревкою схватить за язык его?
JOB|40|26|вденешь ли кольцо в ноздри его? проколешь ли иглою челюсть его?
JOB|40|27|будет ли он много умолять тебя и будет ли говорить с тобою кротко?
JOB|40|28|сделает ли он договор с тобою, и возьмешь ли его навсегда себе в рабы?
JOB|40|29|станешь ли забавляться им, как птичкою, и свяжешь ли его для девочек твоих?
JOB|40|30|будут ли продавать его товарищи ловли, разделят ли его между Хананейскими купцами?
JOB|40|31|можешь ли пронзить кожу его копьем и голову его рыбачьею острогою?
JOB|40|32|Клади на него руку твою, и помни о борьбе: вперед не будешь.
JOB|41|1|Надежда тщетна: не упадешь ли от одного взгляда его?
JOB|41|2|Нет столь отважного, который осмелился бы потревожить его; кто же может устоять перед Моим лицем?
JOB|41|3|Кто предварил Меня, чтобы Мне воздавать ему? под всем небом все Мое.
JOB|41|4|Не умолчу о членах его, о силе и красивой соразмерности их.
JOB|41|5|Кто может открыть верх одежды его, кто подойдет к двойным челюстям его?
JOB|41|6|Кто может отворить двери лица его? круг зубов его – ужас;
JOB|41|7|крепкие щиты его – великолепие; они скреплены как бы твердою печатью;
JOB|41|8|один к другому прикасается близко, так что и воздух не проходит между ними;
JOB|41|9|один с другим лежат плотно, сцепились и не раздвигаются.
JOB|41|10|От его чихания показывается свет; глаза у него как ресницы зари;
JOB|41|11|из пасти его выходят пламенники, выскакивают огненные искры;
JOB|41|12|из ноздрей его выходит дым, как из кипящего горшка или котла.
JOB|41|13|Дыхание его раскаляет угли, и из пасти его выходит пламя.
JOB|41|14|На шее его обитает сила, и перед ним бежит ужас.
JOB|41|15|Мясистые части тела его сплочены между собою твердо, не дрогнут.
JOB|41|16|Сердце его твердо, как камень, и жестко, как нижний жернов.
JOB|41|17|Когда он поднимается, силачи в страхе, совсем теряются от ужаса.
JOB|41|18|Меч, коснувшийся его, не устоит, ни копье, ни дротик, ни латы.
JOB|41|19|Железо он считает за солому, медь – за гнилое дерево.
JOB|41|20|Дочь лука не обратит его в бегство; пращные камни обращаются для него в плеву.
JOB|41|21|Булава считается у него за соломину; свисту дротика он смеется.
JOB|41|22|Под ним острые камни, и он на острых камнях лежит в грязи.
JOB|41|23|Он кипятит пучину, как котел, и море претворяет в кипящую мазь;
JOB|41|24|оставляет за собою светящуюся стезю; бездна кажется сединою.
JOB|41|25|Нет на земле подобного ему; он сотворен бесстрашным;
JOB|41|26|на все высокое смотрит смело; он царь над всеми сынами гордости.
JOB|42|1|И отвечал Иов Господу и сказал:
JOB|42|2|знаю, что Ты все можешь, и что намерение Твое не может быть остановлено.
JOB|42|3|Кто сей, омрачающий Провидение, ничего не разумея? – Так, я говорил о том, чего не разумел, о делах чудных для меня, которых я не знал.
JOB|42|4|Выслушай, [взывал я,] и я буду говорить, и что буду спрашивать у Тебя, объясни мне.
JOB|42|5|Я слышал о Тебе слухом уха; теперь же мои глаза видят Тебя;
JOB|42|6|поэтому я отрекаюсь и раскаиваюсь в прахе и пепле.
JOB|42|7|И было после того, как Господь сказал слова те Иову, сказал Господь Елифазу Феманитянину: горит гнев Мой на тебя и на двух друзей твоих за то, что вы говорили о Мне не так верно, как раб Мой Иов.
JOB|42|8|Итак возьмите себе семь тельцов и семь овнов и пойдите к рабу Моему Иову и принесите за себя жертву; и раб Мой Иов помолится за вас, ибо только лице его Я приму, дабы не отвергнуть вас за то, что вы говорили о Мне не так верно, как раб Мой Иов.
JOB|42|9|И пошли Елифаз Феманитянин и Вилдад Савхеянин и Софар Наамитянин, и сделали так, как Господь повелел им, – и Господь принял лице Иова.
JOB|42|10|И возвратил Господь потерю Иова, когда он помолился за друзей своих; и дал Господь Иову вдвое больше того, что он имел прежде.
JOB|42|11|Тогда пришли к нему все братья его и все сестры его и все прежние знакомые его, и ели с ним хлеб в доме его, и тужили с ним, и утешали его за все зло, которое Господь навел на него, и дали ему каждый по кесите и по золотому кольцу.
JOB|42|12|И благословил Бог последние дни Иова более, нежели прежние: у него было четырнадцать тысяч мелкого скота, шесть тысяч верблюдов, тысяча пар волов и тысяча ослиц.
JOB|42|13|И было у него семь сыновей и три дочери.
JOB|42|14|И нарек он имя первой Емима, имя второй – Кассия, а имя третьей – Керенгаппух.
JOB|42|15|И не было на всей земле таких прекрасных женщин, как дочери Иова, и дал им отец их наследство между братьями их.
JOB|42|16|После того Иов жил сто сорок лет, и видел сыновей своих и сыновей сыновних до четвертого рода;
JOB|42|17|и умер Иов в старости, насыщенный днями.
