JONAH|1|1|耶和华的话临到 亚米太 的儿子 约拿 ，说：
JONAH|1|2|“起来，到 尼尼微 大城去，向其中的居民宣告，因为他们的恶已达到我面前。”
JONAH|1|3|约拿 却起身，逃往 他施 去躲避耶和华。他下到 约帕 ，遇见一条船要往 他施 去。 约拿 付了船费，就上船，与船上的人同往 他施 ，为要躲避耶和华。
JONAH|1|4|耶和华在海上刮起大风，海就狂风大作，船几乎破裂。
JONAH|1|5|水手都惧怕，各人哀求自己的神明。他们把船上的货物抛进海里，为要减轻载重。 约拿 却下到舱底，躺卧沉睡。
JONAH|1|6|船长到他那里，对他说：“你怎么还在沉睡呢？起来，求告你的神明，或者神明顾念我们，使我们不致灭亡。”
JONAH|1|7|船上的人彼此说：“来吧，我们来抽签，看看这灾难临到我们是因谁的缘故。”于是他们就抽签，抽出 约拿 来。
JONAH|1|8|他们对 约拿 说：“请你告诉我们，这灾难临到我们是因谁的缘故呢？你做什么行业？你从哪里来？你是哪一国的人？属哪一族？”
JONAH|1|9|他说：“我是 希伯来 人，我敬畏耶和华，天上的上帝，他创造了沧海和陆地。”
JONAH|1|10|那些人就大大惧怕，对他说：“你做的是什么事呢？”原来他们已经知道他在躲避耶和华，因为他告诉了他们。
JONAH|1|11|海浪越来越汹涌，他们就问他说：“我们当向你做什么，才能使海浪平静呢？”
JONAH|1|12|他对他们说：“你们把我抬起来，抛进海里，海就会平静了；我知道你们遭遇这大风浪是因我的缘故。”
JONAH|1|13|然而那些人竭力划桨，想要把船靠回陆地，却是不能；因风浪愈来愈大，扑向他们。
JONAH|1|14|于是他们求告耶和华说：“耶和华啊，求求你不要因这人的性命使我们灭亡，不要使流无辜人血的罪归给我们；因为你－耶和华随自己的旨意行事。”
JONAH|1|15|他们把 约拿 抬起来，抛进海里，海的狂浪就平息了。
JONAH|1|16|那些人就大大惧怕耶和华，向耶和华献祭许愿。
JONAH|1|17|耶和华安排一条大鱼吞下 约拿 ， 约拿 在鱼腹中三日三夜。
JONAH|2|1|约拿 在鱼腹中向耶和华－他的上帝祷告，
JONAH|2|2|说： “我在患难中求告耶和华， 他就应允我； 我从阴间的深处呼求， 你就俯听我的声音。
JONAH|2|3|你将我投下深渊， 直到海心； 大水环绕我， 你的波浪洪涛漫过我身。
JONAH|2|4|我说：‘我从你眼前被驱逐， 然而我仍要仰望你的圣殿。’
JONAH|2|5|众水环绕我，几乎淹没我； 深渊围住我； 海草缠绕我的头。
JONAH|2|6|我下沉到山的根基， 地的门闩将我永远关住。 耶和华－我的上帝啊， 你却将我的性命从地府里救出来。
JONAH|2|7|我心灵发昏时， 就想起耶和华。 我的祷告进入你的圣殿， 达到你面前。
JONAH|2|8|那信奉虚无神明 的人， 丢弃自己的慈爱；
JONAH|2|9|但我要以感谢的声音向你献祭。 我所许的愿，我必偿还。 救恩出于耶和华。”
JONAH|2|10|耶和华吩咐那鱼，鱼就把 约拿 吐在陆地上。
JONAH|3|1|耶和华的话第二次临到 约拿 ，说：
JONAH|3|2|“起来，到 尼尼微 大城去，把我告诉你的信息向其中的居民宣告。”
JONAH|3|3|约拿 就照耶和华的话起来，到 尼尼微 去。 尼尼微 是一座极大的城，约有三天的路程。
JONAH|3|4|约拿 进城，走了一天，宣告说：“再过四十天， 尼尼微 要倾覆了！”
JONAH|3|5|尼尼微 人就信服上帝，宣告禁食，从最大的到最小的都穿上麻衣。
JONAH|3|6|这消息传到 尼尼微 王那里，他就从宝座起来，脱下朝服，披上麻布，坐在灰中。
JONAH|3|7|他叫人通告 尼尼微 全城，说：“王和大臣有令，人、畜、牛、羊都不可尝任何东西，不可吃，也不可喝水。
JONAH|3|8|人与牲畜都要披上麻布，切切求告上帝。各人要回转离开恶道，离弃自己掌中的残暴。
JONAH|3|9|谁知道上帝也许会回心转意，不发烈怒，使我们不致灭亡。”
JONAH|3|10|上帝察看他们的行为，见他们离开恶道，上帝就改变心意，原先所说要降与他们的灾难，他不降了。
JONAH|4|1|这事令 约拿 大大不悦，甚至发怒。
JONAH|4|2|他就向耶和华祷告，说：“耶和华啊，这不就是我仍在本国的时候所说的吗？我知道你是有恩惠，有怜悯的上帝，不轻易发怒，有丰盛的慈爱，并且会改变心意，不降那灾难。我就是因为这样，才急速逃往 他施 去的呀！
JONAH|4|3|耶和华啊，现在求你取走我的性命吧！因为我死了比活着更好。”
JONAH|4|4|耶和华说：“你这样发怒，对吗？”
JONAH|4|5|约拿 出城，坐在城的东边，在那里为自己搭了一座棚。他坐在棚子的荫下，要看看城里会发生什么事。
JONAH|4|6|耶和华上帝安排了一棵蓖麻，使它生长高过 约拿 ，影子遮盖他的头，使他免受苦难； 约拿 因这棵蓖麻大大欢喜。
JONAH|4|7|次日黎明，上帝却安排一条虫来咬这蓖麻，以致枯干。
JONAH|4|8|太阳出来的时候，上帝安排炎热的东风，太阳曝晒 约拿 的头，使他发昏，他就为自己求死，说：“我死了比活着更好！”
JONAH|4|9|上帝对 约拿 说：“你因这棵蓖麻这样发怒，对吗？”他说：“我发怒以至于死，都是对的！”
JONAH|4|10|耶和华说：“这棵蓖麻你没有为它操劳，也不是你使它长大的；它一夜生长，一夜枯死，你尚且爱惜；
JONAH|4|11|何况这 尼尼微 大城，其中不能分辨左右手的就有十二万多人，还有许多牲畜，我岂能不爱惜呢？”
