NUM|1|1|The LORD spoke to Moses in the wilderness of Sinai, in the tent of meeting, on the first day of the second month, in the second year after they had come out of the land of Egypt, saying,
NUM|1|2|"Take a census of all the congregation of the people of Israel, by clans, by fathers' houses, according to the number of names, every male, head by head.
NUM|1|3|From twenty years old and upward, all in Israel who are able to go to war, you and Aaron shall list them, company by company.
NUM|1|4|And there shall be with you a man from each tribe, each man being the head of the house of his fathers.
NUM|1|5|And these are the names of the men who shall assist you. From Reuben, Elizur the son of Shedeur;
NUM|1|6|from Simeon, Shelumiel the son of Zurishaddai;
NUM|1|7|from Judah, Nahshon the son of Amminadab;
NUM|1|8|from Issachar, Nethanel the son of Zuar;
NUM|1|9|from Zebulun, Eliab the son of Helon;
NUM|1|10|from the sons of Joseph, from Ephraim, Elishama the son of Ammihud, and from Manasseh, Gamaliel the son of Pedahzur;
NUM|1|11|from Benjamin, Abidan the son of Gideoni;
NUM|1|12|from Dan, Ahiezer the son of Ammishaddai;
NUM|1|13|from Asher, Pagiel the son of Ochran;
NUM|1|14|from Gad, Eliasaph the son of Deuel;
NUM|1|15|from Naphtali, Ahira the son of Enan."
NUM|1|16|These were the ones chosen from the congregation, the chiefs of their ancestral tribes, the heads of the clans of Israel.
NUM|1|17|Moses and Aaron took these men who had been named,
NUM|1|18|and on the first day of the second month, they assembled the whole congregation together, who registered themselves by clans, by fathers' houses, according to the number of names from twenty years old and upward, head by head,
NUM|1|19|as the LORD commanded Moses. So he listed them in the wilderness of Sinai.
NUM|1|20|The people of Reuben, Israel's firstborn, their generations, by their clans, by their fathers' houses, according to the number of names, head by head, every male from twenty years old and upward, all who were able to go to war:
NUM|1|21|those listed of the tribe of Reuben were 46,500.
NUM|1|22|Of the people of Simeon, their generations, by their clans, by their fathers' houses, those of them who were listed, according to the number of names, head by head, every male from twenty years old and upward, all who were able to go to war:
NUM|1|23|those listed of the tribe of Simeon were 59,300.
NUM|1|24|Of the people of Gad, their generations, by their clans, by their fathers' houses, according to the number of the names, from twenty years old and upward, all who were able to go to war:
NUM|1|25|those listed of the tribe of Gad were 45,650.
NUM|1|26|Of the people of Judah, their generations, by their clans, by their fathers' houses, according to the number of names, from twenty years old and upward, every man able to go to war:
NUM|1|27|those listed of the tribe of Judah were 74,600.
NUM|1|28|Of the people of Issachar, their generations, by their clans, by their fathers' houses, according to the number of names, from twenty years old and upward, every man able to go to war:
NUM|1|29|those listed of the tribe of Issachar were 54,400.
NUM|1|30|Of the people of Zebulun, their generations, by their clans, by their fathers' houses, according to the number of names, from twenty years old and upward, every man able to go to war:
NUM|1|31|those listed of the tribe of Zebulun were 57,400.
NUM|1|32|Of the people of Joseph, namely, of the people of Ephraim, their generations, by their clans, by their fathers' houses, according to the number of names, from twenty years old and upward, every man able to go to war:
NUM|1|33|those listed of the tribe of Ephraim were 40,500.
NUM|1|34|Of the people of Manasseh, their generations, by their clans, by their fathers' houses, according to the number of names, from twenty years old and upward, every man able to go to war:
NUM|1|35|those listed of the tribe of Manasseh were 32,200.
NUM|1|36|Of the people of Benjamin, their generations, by their clans, by their fathers' houses, according to the number of names, from twenty years old and upward, every man able to go to war:
NUM|1|37|those listed of the tribe of Benjamin were 35,400.
NUM|1|38|Of the people of Dan, their generations, by their clans, by their fathers' houses, according to the number of names, from twenty years old and upward, every man able to go to war:
NUM|1|39|those listed of the tribe of Dan were 62,700.
NUM|1|40|Of the people of Asher, their generations, by their clans, by their fathers' houses, according to the number of names, from twenty years old and upward, every man able to go to war:
NUM|1|41|those listed of the tribe of Asher were 41,500.
NUM|1|42|Of the people of Naphtali, their generations, by their clans, by their fathers' houses, according to the number of names, from twenty years old and upward, every man able to go to war:
NUM|1|43|those listed of the tribe of Naphtali were 53,400.
NUM|1|44|These are those who were listed, whom Moses and Aaron listed with the help of the chiefs of Israel, twelve men, each representing his fathers' house.
NUM|1|45|So all those listed of the people of Israel, by their fathers' houses, from twenty years old and upward, every man able to go to war in Israel-
NUM|1|46|all those listed were 603,550.
NUM|1|47|But the Levites were not listed along with them by their ancestral tribe.
NUM|1|48|For the LORD spoke to Moses, saying,
NUM|1|49|"Only the tribe of Levi you shall not list, and you shall not take a census of them among the people of Israel.
NUM|1|50|But appoint the Levites over the tabernacle of the testimony, and over all its furnishings, and over all that belongs to it. They are to carry the tabernacle and all its furnishings, and they shall take care of it and shall camp around the tabernacle.
NUM|1|51|When the tabernacle is to set out, the Levites shall take it down, and when the tabernacle is to be pitched, the Levites shall set it up. And if any outsider comes near, he shall be put to death.
NUM|1|52|The people of Israel shall pitch their tents by their companies, each man in his own camp and each man by his own standard.
NUM|1|53|But the Levites shall camp around the tabernacle of the testimony, so that there may be no wrath on the congregation of the people of Israel. And the Levites shall keep guard over the tabernacle of the testimony."
NUM|1|54|Thus did the people of Israel; they did according to all that the LORD commanded Moses.
NUM|2|1|The LORD spoke to Moses and Aaron, saying,
NUM|2|2|"The people of Israel shall camp each by his own standard, with the banners of their fathers' houses. They shall camp facing the tent of meeting on every side.
NUM|2|3|Those to camp on the east side toward the sunrise shall be of the standard of the camp of Judah by their companies, the chief of the people of Judah being Nahshon the son of Amminadab,
NUM|2|4|his company as listed being 74,600.
NUM|2|5|Those to camp next to him shall be the tribe of Issachar, the chief of the people of Issachar being Nethanel the son of Zuar,
NUM|2|6|his company as listed being 54,400.
NUM|2|7|Then the tribe of Zebulun, the chief of the people of Zebulun being Eliab the son of Helon,
NUM|2|8|his company as listed being 57,400.
NUM|2|9|All those listed of the camp of Judah, by their companies, were 186,400. They shall set out first on the march.
NUM|2|10|"On the south side shall be the standard of the camp of Reuben by their companies, the chief of the people of Reuben being Elizur the son of Shedeur,
NUM|2|11|his company as listed being 46,500.
NUM|2|12|And those to camp next to him shall be the tribe of Simeon, the chief of the people of Simeon being Shelumiel the son of Zurishaddai,
NUM|2|13|his company as listed being 59,300.
NUM|2|14|Then the tribe of Gad, the chief of the people of Gad being Eliasaph the son of Reuel,
NUM|2|15|his company as listed being 45,650.
NUM|2|16|All those listed of the camp of Reuben, by their companies, were 151,450. They shall set out second.
NUM|2|17|"Then the tent of meeting shall set out, with the camp of the Levites in the midst of the camps; as they camp, so shall they set out, each in position, standard by standard.
NUM|2|18|"On the west side shall be the standard of the camp of Ephraim by their companies, the chief of the people of Ephraim being Elishama the son of Ammihud,
NUM|2|19|his company as listed being 40,500.
NUM|2|20|And next to him shall be the tribe of Manasseh, the chief of the people of Manasseh being Gamaliel the son of Pedahzur,
NUM|2|21|his company as listed being 32,200.
NUM|2|22|Then the tribe of Benjamin, the chief of the people of Benjamin being Abidan the son of Gideoni,
NUM|2|23|his company as listed being 35,400.
NUM|2|24|All those listed of the camp of Ephraim, by their companies, were 108,100. They shall set out third on the march.
NUM|2|25|"On the north side shall be the standard of the camp of Dan by their companies, the chief of the people of Dan being Ahiezer the son of Ammishaddai,
NUM|2|26|his company as listed being 62,700.
NUM|2|27|And those to camp next to him shall be the tribe of Asher, the chief of the people of Asher being Pagiel the son of Ochran,
NUM|2|28|his company as listed being 41,500.
NUM|2|29|Then the tribe of Naphtali, the chief of the people of Naphtali being Ahira the son of Enan,
NUM|2|30|his company as listed being 53,400.
NUM|2|31|All those listed of the camp of Dan were 157,600. They shall set out last, standard by standard."
NUM|2|32|These are the people of Israel as listed by their fathers' houses. All those listed in the camps by their companies were 603,550.
NUM|2|33|But the Levites were not listed among the people of Israel, as the LORD commanded Moses.
NUM|2|34|Thus did the people of Israel. According to all that the LORD commanded Moses, so they camped by their standards, and so they set out, each one in his clan, according to his fathers' house.
NUM|3|1|These are the generations of Aaron and Moses at the time when the LORD spoke with Moses on Mount Sinai.
NUM|3|2|These are the names of the sons of Aaron: Nadab the firstborn, and Abihu, Eleazar, and Ithamar.
NUM|3|3|These are the names of the sons of Aaron, the anointed priests, whom he ordained to serve as priests.
NUM|3|4|But Nadab and Abihu died before the LORD when they offered unauthorized fire before the LORD in the wilderness of Sinai, and they had no children. So Eleazar and Ithamar served as priests in the lifetime of Aaron their father.
NUM|3|5|And the LORD spoke to Moses, saying,
NUM|3|6|"Bring the tribe of Levi near, and set them before Aaron the priest, that they may minister to him.
NUM|3|7|They shall keep guard over him and over the whole congregation before the tent of meeting, as they minister at the tabernacle.
NUM|3|8|They shall guard all the furnishings of the tent of meeting, and keep guard over the people of Israel as they minister at the tabernacle.
NUM|3|9|And you shall give the Levites to Aaron and his sons; they are wholly given to him from among the people of Israel.
NUM|3|10|And you shall appoint Aaron and his sons, and they shall guard their priesthood. But if any outsider comes near, he shall be put to death."
NUM|3|11|And the LORD spoke to Moses, saying,
NUM|3|12|"Behold, I have taken the Levites from among the people of Israel instead of every firstborn who opens the womb among the people of Israel. The Levites shall be mine,
NUM|3|13|for all the firstborn are mine. On the day that I struck down all the firstborn in the land of Egypt, I consecrated for my own all the firstborn in Israel, both of man and of beast. They shall be mine: I am the LORD."
NUM|3|14|And the LORD spoke to Moses in the wilderness of Sinai, saying,
NUM|3|15|"List the sons of Levi, by fathers' houses and by clans; every male from a month old and upward you shall list."
NUM|3|16|So Moses listed them according to the word of the LORD, as he was commanded.
NUM|3|17|And these were the sons of Levi by their names: Gershon and Kohath and Merari.
NUM|3|18|And these are the names of the sons of Gershon by their clans: Libni and Shimei.
NUM|3|19|And the sons of Kohath by their clans: Amram, Izhar, Hebron, and Uzziel.
NUM|3|20|And the sons of Merari by their clans: Mahli and Mushi. These are the clans of the Levites, by their fathers' houses.
NUM|3|21|To Gershon belonged the clan of the Libnites and the clan of the Shimeites; these were the clans of the Gershonites.
NUM|3|22|Their listing according to the number of all the males from a month old and upward was 7,500.
NUM|3|23|The clans of the Gershonites were to camp behind the tabernacle on the west,
NUM|3|24|with Eliasaph, the son of Lael as chief of the fathers' house of the Gershonites.
NUM|3|25|And the guard duty of the sons of Gershon in the tent of meeting involved the tabernacle, the tent with its covering, the screen for the entrance of the tent of meeting,
NUM|3|26|the hangings of the court, the screen for the door of the court that is around the tabernacle and the altar, and its cords- all the service connected with these.
NUM|3|27|To Kohath belonged the clan of the Amramites and the clan of the Izharites and the clan of the Hebronites and the clan of the Uzzielites; these are the clans of the Kohathites.
NUM|3|28|According to the number of all the males, from a month old and upward, there were 8,600, keeping guard over the sanctuary.
NUM|3|29|The clans of the sons of Kohath were to camp on the south side of the tabernacle,
NUM|3|30|with Elizaphan the son of Uzziel as chief of the fathers' house of the clans of the Kohathites.
NUM|3|31|And their guard duty involved the ark, the table, the lampstand, the altars, the vessels of the sanctuary with which the priests minister, and the screen; all the service connected with these.
NUM|3|32|And Eleazar the son of Aaron the priest was to be chief over the chiefs of the Levites, and to have oversight of those who kept guard over the sanctuary.
NUM|3|33|To Merari belonged the clan of the Mahlites and the clan of the Mushites: these are the clans of Merari.
NUM|3|34|Their listing according to the number of all the males from a month old and upward was 6,200.
NUM|3|35|And the chief of the fathers' house of the clans of Merari was Zuriel the son of Abihail. They were to camp on the north side of the tabernacle.
NUM|3|36|And the appointed guard duty of the sons of Merari involved the frames of the tabernacle, the bars, the pillars, the bases, and all their accessories; all the service connected with these;
NUM|3|37|also the pillars around the court, with their bases and pegs and cords.
NUM|3|38|Those who were to camp before the tabernacle on the east, before the tent of meeting toward the sunrise, were Moses and Aaron and his sons, guarding the sanctuary itself, to protect the people of Israel. And any outsider who came near was to be put to death.
NUM|3|39|All those listed among the Levites, whom Moses and Aaron listed at the commandment of the LORD, by clans, all the males from a month old and upward, were 22,000.
NUM|3|40|And the LORD said to Moses, "List all the firstborn males of the people of Israel, from a month old and upward, taking the number of their names.
NUM|3|41|And you shall take the Levites for me- I am the LORD- instead of all the firstborn among the people of Israel, and the cattle of the Levites instead of all the firstborn among the cattle of the people of Israel."
NUM|3|42|So Moses listed all the firstborn among the people of Israel, as the LORD commanded him.
NUM|3|43|And all the firstborn males, according to the number of names, from a month old and upward as listed were 22,273.
NUM|3|44|And the LORD spoke to Moses, saying,
NUM|3|45|"Take the Levites instead of all the firstborn among the people of Israel, and the cattle of the Levites instead of their cattle. The Levites shall be mine: I am the LORD.
NUM|3|46|And as the redemption price for the 273 of the firstborn of the people of Israel, over and above the number of the male Levites,
NUM|3|47|you shall take five shekels per head; you shall take them according to the shekel of the sanctuary (the shekel of twenty gerahs),
NUM|3|48|and give the money to Aaron and his sons as the redemption price for those who are over."
NUM|3|49|So Moses took the redemption money from those who were over and above those redeemed by the Levites.
NUM|3|50|From the firstborn of the people of Israel he took the money, 1,365 shekels, by the shekel of the sanctuary.
NUM|3|51|And Moses gave the redemption money to Aaron and his sons, according to the word of the LORD, as the LORD commanded Moses.
NUM|4|1|The LORD spoke to Moses and Aaron, saying,
NUM|4|2|"Take a census of the sons of Kohath from among the sons of Levi, by their clans and their fathers' houses,
NUM|4|3|from thirty years old up to fifty years old, all who can come on duty, to do the work in the tent of meeting.
NUM|4|4|This is the service of the sons of Kohath in the tent of meeting: the most holy things.
NUM|4|5|When the camp is to set out, Aaron and his sons shall go in and take down the veil of the screen and cover the ark of the testimony with it.
NUM|4|6|Then they shall put on it a covering of goatskin and spread on top of that a cloth all of blue, and shall put in its poles.
NUM|4|7|And over the table of the bread of the Presence they shall spread a cloth of blue and put on it the plates, the dishes for incense, the bowls, and the flagons for the drink offering; the regular show bread also shall be on it.
NUM|4|8|Then they shall spread over them a cloth of scarlet and cover the same with a covering of goatskin, and shall put in its poles.
NUM|4|9|And they shall take a cloth of blue and cover the lampstand for the light, with its lamps, its tongs, its trays, and all the vessels for oil with which it is supplied.
NUM|4|10|And they shall put it with all its utensils in a covering of goatskin and put it on the carrying frame.
NUM|4|11|And over the golden altar they shall spread a cloth of blue and cover it with a covering of goatskin, and shall put in its poles.
NUM|4|12|And they shall take all the vessels of the service that are used in the sanctuary and put them in a cloth of blue and cover them with a covering of goatskin and put them on the carrying frame.
NUM|4|13|And they shall take away the ashes from the altar and spread a purple cloth over it.
NUM|4|14|And they shall put on it all the utensils of the altar, which are used for the service there, the fire pans, the forks, the shovels, and the basins, all the utensils of the altar; and they shall spread on it a covering of goatskin, and shall put in its poles.
NUM|4|15|And when Aaron and his sons have finished covering the sanctuary and all the furnishings of the sanctuary, as the camp sets out, after that the sons of Kohath shall come to carry these, but they must not touch the holy things, lest they die. These are the things of the tent of meeting that the sons of Kohath are to carry.
NUM|4|16|"And Eleazar the son of Aaron the priest shall have charge of the oil for the light, the fragrant incense, the regular grain offering, and the anointing oil, with the oversight of the whole tabernacle and all that is in it, of the sanctuary and its vessels."
NUM|4|17|The LORD spoke to Moses and Aaron, saying,
NUM|4|18|"Let not the tribe of the clans of the Kohathites be destroyed from among the Levites,
NUM|4|19|but deal thus with them, that they may live and not die when they come near to the most holy things: Aaron and his sons shall go in and appoint them each to his task and to his burden,
NUM|4|20|but they shall not go in to look on the holy things even for a moment, lest they die."
NUM|4|21|The LORD spoke to Moses, saying,
NUM|4|22|"Take a census of the sons of Gershon also, by their fathers' houses and by their clans.
NUM|4|23|From thirty years old up to fifty years old, you shall list them, all who can come to do duty, to do service in the tent of meeting.
NUM|4|24|This is the service of the clans of the Gershonites, in serving and bearing burdens:
NUM|4|25|they shall carry the curtains of the tabernacle and the tent of meeting with its covering and the covering of goatskin that is on top of it and the screen for the entrance of the tent of meeting
NUM|4|26|and the hangings of the court and the screen for the entrance of the gate of the court that is around the tabernacle and the altar, and their cords and all the equipment for their service. And they shall do all that needs to be done with regard to them.
NUM|4|27|All the service of the sons of the Gershonites shall be at the command of Aaron and his sons, in all that they are to carry and in all that they have to do. And you shall assign to their charge all that they are to carry.
NUM|4|28|This is the service of the clans of the sons of the Gershonites in the tent of meeting, and their guard duty is to be under the direction of Ithamar the son of Aaron the priest.
NUM|4|29|"As for the sons of Merari, you shall list them by their clans and their fathers' houses.
NUM|4|30|From thirty years old up to fifty years old, you shall list them, everyone who can come on duty, to do the service of the tent of meeting.
NUM|4|31|And this is what they are charged to carry, as the whole of their service in the tent of meeting: the frames of the tabernacle, with its bars, pillars, and bases,
NUM|4|32|and the pillars around the court with their bases, pegs, and cords, with all their equipment and all their accessories. And you shall list by name the objects that they are required to carry.
NUM|4|33|This is the service of the clans of the sons of Merari, the whole of their service in the tent of meeting, under the direction of Ithamar the son of Aaron the priest."
NUM|4|34|And Moses and Aaron and the chiefs of the congregation listed the sons of the Kohathites, by their clans and their fathers' houses,
NUM|4|35|from thirty years old up to fifty years old, everyone who could come on duty, for service in the tent of meeting;
NUM|4|36|and those listed by clans were 2,750.
NUM|4|37|This was the list of the clans of the Kohathites, all who served in the tent of meeting, whom Moses and Aaron listed according to the commandment of the LORD by Moses.
NUM|4|38|Those listed of the sons of Gershon, by their clans and their fathers' houses,
NUM|4|39|from thirty years old up to fifty years old, everyone who could come on duty for service in the tent of meeting-
NUM|4|40|those listed by their clans and their fathers' houses were 2,630.
NUM|4|41|This was the list of the clans of the sons of Gershon, all who served in the tent of meeting, whom Moses and Aaron listed according to the commandment of the LORD.
NUM|4|42|Those listed of the clans of the sons of Merari, by their clans and their fathers' houses,
NUM|4|43|from thirty years old up to fifty years old, everyone who could come on duty, for service in the tent of meeting-
NUM|4|44|those listed by clans were 3,200.
NUM|4|45|This was the list of the clans of the sons of Merari, whom Moses and Aaron listed according to the commandment of the LORD by Moses.
NUM|4|46|All those who were listed of the Levites, whom Moses and Aaron and the chiefs of Israel listed, by their clans and their fathers' houses,
NUM|4|47|from thirty years old up to fifty years old, everyone who could come to do the service of ministry and the service of bearing burdens in the tent of meeting,
NUM|4|48|those listed were 8,580.
NUM|4|49|According to the commandment of the LORD through Moses they were listed, each one with his task of serving or carrying. Thus they were listed by him, as the LORD commanded Moses.
NUM|5|1|The LORD spoke to Moses, saying,
NUM|5|2|"Command the people of Israel that they put out of the camp everyone who is leprous or has a discharge and everyone who is unclean through contact with the dead.
NUM|5|3|You shall put out both male and female, putting them outside the camp, that they may not defile their camp, in the midst of which I dwell."
NUM|5|4|And the people of Israel did so, and put them outside the camp; as the LORD said to Moses, so the people of Israel did.
NUM|5|5|And the LORD spoke to Moses, saying,
NUM|5|6|"Speak to the people of Israel, When a man or woman commits any of the sins that people commit by breaking faith with the LORD, and that person realizes his guilt,
NUM|5|7|he shall confess his sin that he has committed. And he shall make full restitution for his wrong, adding a fifth to it and giving it to him to whom he did the wrong.
NUM|5|8|But if the man has no next of kin to whom restitution may be made for the wrong, the restitution for wrong shall go to the LORD for the priest, in addition to the ram of atonement with which atonement is made for him.
NUM|5|9|And every contribution, all the holy donations of the people of Israel, which they bring to the priest, shall be his.
NUM|5|10|Each one shall keep his holy donations: whatever anyone gives to the priest shall be his."
NUM|5|11|And the LORD spoke to Moses, saying,
NUM|5|12|"Speak to the people of Israel, If any man's wife goes astray and breaks faith with him,
NUM|5|13|if a man lies with her sexually, and it is hidden from the eyes of her husband, and she is undetected though she has defiled herself, and there is no witness against her, since she was not taken in the act,
NUM|5|14|and if the spirit of jealousy comes over him and he is jealous of his wife who has defiled herself, or if the spirit of jealousy comes over him and he is jealous of his wife, though she has not defiled herself,
NUM|5|15|then the man shall bring his wife to the priest and bring the offering required of her, a tenth of an ephah of barley flour. He shall pour no oil on it and put no frankincense on it, for it is a grain offering of jealousy, a grain offering of remembrance, bringing iniquity to remembrance.
NUM|5|16|"And the priest shall bring her near and set her before the LORD.
NUM|5|17|And the priest shall take holy water in an earthenware vessel and take some of the dust that is on the floor of the tabernacle and put it into the water.
NUM|5|18|And the priest shall set the woman before the LORD and unbind the hair of the woman's head and place in her hands the grain offering of remembrance, which is the grain offering of jealousy. And in his hand the priest shall have the water of bitterness that brings the curse.
NUM|5|19|Then the priest shall make her take an oath, saying, 'If no man has lain with you, and if you have not turned aside to uncleanness while you were under your husband's authority, be free from this water of bitterness that brings the curse.
NUM|5|20|But if you have gone astray, though you are under your husband's authority, and if you have defiled yourself, and some man other than your husband has lain with you,
NUM|5|21|then' (let the priest make the woman take the oath of the curse, and say to the woman) 'the LORD make you a curse and an oath among your people, when the LORD makes your thigh fall away and your body swell.
NUM|5|22|May this water that brings the curse pass into your bowels and make your womb swell and your thigh fall away.' And the woman shall say, 'Amen, Amen.'
NUM|5|23|"Then the priest shall write these curses in a book and wash them off into the water of bitterness.
NUM|5|24|And he shall make the woman drink the water of bitterness that brings the curse, and the water that brings the curse shall enter into her and cause bitter pain.
NUM|5|25|And the priest shall take the grain offering of jealousy out of the woman's hand and shall wave the grain offering before the LORD and bring it to the altar.
NUM|5|26|And the priest shall take a handful of the grain offering, as its memorial portion, and burn it on the altar, and afterward shall make the woman drink the water.
NUM|5|27|And when he has made her drink the water, then, if she has defiled herself and has broken faith with her husband, the water that brings the curse shall enter into her and cause bitter pain, and her womb shall swell, and her thigh shall fall away, and the woman shall become a curse among her people.
NUM|5|28|But if the woman has not defiled herself and is clean, then she shall be free and shall conceive children.
NUM|5|29|"This is the law in cases of jealousy, when a wife, though under her husband's authority, goes astray and defiles herself,
NUM|5|30|or when the spirit of jealousy comes over a man and he is jealous of his wife. Then he shall set the woman before the LORD, and the priest shall carry out for her all this law.
NUM|5|31|The man shall be free from iniquity, but the woman shall bear her iniquity."
NUM|6|1|And the LORD spoke to Moses, saying,
NUM|6|2|"Speak to the people of Israel and say to them, When either a man or a woman makes a special vow, the vow of a Nazirite, to separate himself to the LORD,
NUM|6|3|he shall separate himself from wine and strong drink. He shall drink no vinegar made from wine or strong drink and shall not drink any juice of grapes or eat grapes, fresh or dried.
NUM|6|4|All the days of his separation he shall eat nothing that is produced by the grapevine, not even the seeds or the skins.
NUM|6|5|"All the days of his vow of separation, no razor shall touch his head. Until the time is completed for which he separates himself to the LORD, he shall be holy. He shall let the locks of hair of his head grow long.
NUM|6|6|"All the days that he separates himself to the LORD he shall not go near a dead body.
NUM|6|7|Not even for his father or for his mother, for brother or sister, if they die, shall he make himself unclean, because his separation to God is on his head.
NUM|6|8|All the days of his separation he is holy to the LORD.
NUM|6|9|"And if any man dies very suddenly beside him and he defiles his consecrated head, then he shall shave his head on the day of his cleansing; on the seventh day he shall shave it.
NUM|6|10|On the eighth day he shall bring two turtledoves or two pigeons to the priest to the entrance of the tent of meeting,
NUM|6|11|and the priest shall offer one for a sin offering and the other for a burnt offering, and make atonement for him, because he sinned by reason of the dead body. And he shall consecrate his head that same day
NUM|6|12|and separate himself to the LORD for the days of his separation and bring a male lamb a year old for a guilt offering. But the previous period shall be void, because his separation was defiled.
NUM|6|13|"And this is the law for the Nazirite, when the time of his separation has been completed: he shall be brought to the entrance of the tent of meeting,
NUM|6|14|and he shall bring his gift to the LORD, one male lamb a year old without blemish for a burnt offering, and one ewe lamb a year old without blemish as a sin offering, and one ram without blemish as a peace offering,
NUM|6|15|and a basket of unleavened bread, loaves of fine flour mixed with oil, and unleavened wafers smeared with oil, and their grain offering and their drink offerings.
NUM|6|16|And the priest shall bring them before the LORD and offer his sin offering and his burnt offering,
NUM|6|17|and he shall offer the ram as a sacrifice of peace offering to the LORD, with the basket of unleavened bread. The priest shall offer also its grain offering and its drink offering.
NUM|6|18|And the Nazirite shall shave his consecrated head at the entrance of the tent of meeting and shall take the hair from his consecrated head and put it on the fire that is under the sacrifice of the peace offering.
NUM|6|19|And the priest shall take the shoulder of the ram, when it is boiled, and one unleavened loaf out of the basket and one unleavened wafer, and shall put them on the hands of the Nazirite, after he has shaved the hair of his consecration,
NUM|6|20|and the priest shall wave them for a wave offering before the LORD. They are a holy portion for the priest, together with the breast that is waved and the thigh that is contributed. And after that the Nazirite may drink wine.
NUM|6|21|"This is the law of the Nazirite. But if he vows an offering to the LORD above his Nazirite vow, as he can afford, in exact accordance with the vow that he takes, then he shall do in addition to the law of the Nazirite."
NUM|6|22|The LORD spoke to Moses, saying,
NUM|6|23|"Speak to Aaron and his sons, saying, Thus you shall bless the people of Israel: you shall say to them,
NUM|6|24|The LORD bless you and keep you;
NUM|6|25|the LORD make his face to shine upon you and be gracious to you;
NUM|6|26|the LORD lift up his countenance upon you and give you peace.
NUM|6|27|"So shall they put my name upon the people of Israel, and I will bless them."
NUM|7|1|On the day when Moses had finished setting up the tabernacle and had anointed and consecrated it with all its furnishings and had anointed and consecrated the altar with all its utensils,
NUM|7|2|the chiefs of Israel, heads of their fathers' houses, who were the chiefs of the tribes, who were over those who were listed, approached
NUM|7|3|and brought their offerings before the LORD, six wagons and twelve oxen, a wagon for every two of the chiefs, and for each one an ox. They brought them before the tabernacle.
NUM|7|4|Then the LORD said to Moses,
NUM|7|5|"Accept these from them, that they may be used in the service of the tent of meeting, and give them to the Levites, to each man according to his service."
NUM|7|6|So Moses took the wagons and the oxen and gave them to the Levites.
NUM|7|7|Two wagons and four oxen he gave to the sons of Gershon, according to their service.
NUM|7|8|And four wagons and eight oxen he gave to the sons of Merari, according to their service, under the direction of Ithamar the son of Aaron the priest.
NUM|7|9|But to the sons of Kohath he gave none, because they were charged with the service of the holy things that had to be carried on the shoulder.
NUM|7|10|And the chiefs offered offerings for the dedication of the altar on the day it was anointed; and the chiefs offered their offering before the altar.
NUM|7|11|And the LORD said to Moses, "They shall offer their offerings, one chief each day, for the dedication of the altar."
NUM|7|12|He who offered his offering the first day was Nahshon the son of Amminadab, of the tribe of Judah.
NUM|7|13|And his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|14|one golden dish of 10 shekels, full of incense;
NUM|7|15|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|16|one male goat for a sin offering;
NUM|7|17|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Nahshon the son of Amminadab.
NUM|7|18|On the second day Nethanel the son of Zuar, the chief of Issachar, made an offering.
NUM|7|19|He offered for his offering one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|20|one golden dish of 10 shekels, full of incense;
NUM|7|21|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|22|one male goat for a sin offering;
NUM|7|23|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Nethanel the son of Zuar.
NUM|7|24|On the third day Eliab the son of Helon, the chief of the people of Zebulun:
NUM|7|25|his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|26|one golden dish of 10 shekels, full of incense;
NUM|7|27|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|28|one male goat for a sin offering;
NUM|7|29|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Eliab the son of Helon.
NUM|7|30|On the fourth day Elizur the son of Shedeur, the chief of the people of Reuben:
NUM|7|31|his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|32|one golden dish of 10 shekels, full of incense;
NUM|7|33|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|34|one male goat for a sin offering;
NUM|7|35|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Elizur the son of Shedeur.
NUM|7|36|On the fifth day Shelumiel the son of Zurishaddai, the chief of the people of Simeon:
NUM|7|37|his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|38|one golden dish of 10 shekels, full of incense;
NUM|7|39|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|40|one male goat for a sin offering;
NUM|7|41|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Shelumiel the son of Zurishaddai.
NUM|7|42|On the sixth day Eliasaph the son of Deuel, the chief of the people of Gad:
NUM|7|43|his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|44|one golden dish of 10 shekels, full of incense;
NUM|7|45|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|46|one male goat for a sin offering;
NUM|7|47|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Eliasaph the son of Deuel.
NUM|7|48|On the seventh day Elishama the son of Ammihud, the chief of the people of Ephraim:
NUM|7|49|his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|50|one golden dish of 10 shekels, full of incense;
NUM|7|51|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|52|one male goat for a sin offering;
NUM|7|53|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Elishama the son of Ammihud.
NUM|7|54|On the eighth day Gamaliel the son of Pedahzur, the chief of the people of Manasseh:
NUM|7|55|his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|56|one golden dish of 10 shekels, full of incense;
NUM|7|57|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|58|one male goat for a sin offering;
NUM|7|59|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Gamaliel the son of Pedahzur.
NUM|7|60|On the ninth day Abidan the son of Gideoni, the chief of the people of Benjamin:
NUM|7|61|his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|62|one golden dish of 10 shekels, full of incense;
NUM|7|63|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|64|one male goat for a sin offering;
NUM|7|65|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Abidan the son of Gideoni.
NUM|7|66|On the tenth day Ahiezer the son of Ammishaddai, the chief of the people of Dan:
NUM|7|67|his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|68|one golden dish of 10 shekels, full of incense;
NUM|7|69|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|70|one male goat for a sin offering;
NUM|7|71|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Ahiezer the son of Ammishaddai.
NUM|7|72|On the eleventh day Pagiel the son of Ochran, the chief of the people of Asher:
NUM|7|73|his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|74|one golden dish of 10 shekels, full of incense;
NUM|7|75|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|76|one male goat for a sin offering;
NUM|7|77|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Pagiel the son of Ochran.
NUM|7|78|On the twelfth day Ahira the son of Enan, the chief of the people of Naphtali:
NUM|7|79|his offering was one silver plate whose weight was 130 shekels, one silver basin of 70 shekels, according to the shekel of the sanctuary, both of them full of fine flour mixed with oil for a grain offering;
NUM|7|80|one golden dish of 10 shekels, full of incense;
NUM|7|81|one bull from the herd, one ram, one male lamb a year old, for a burnt offering;
NUM|7|82|one male goat for a sin offering;
NUM|7|83|and for the sacrifice of peace offerings, two oxen, five rams, five male goats, and five male lambs a year old. This was the offering of Ahira the son of Enan.
NUM|7|84|This was the dedication offering for the altar on the day when it was anointed, from the chiefs of Israel: twelve silver plates, twelve silver basins, twelve golden dishes,
NUM|7|85|each silver plate weighing 130 shekels and each basin 70, all the silver of the vessels 2,400 shekels according to the shekel of the sanctuary,
NUM|7|86|the twelve golden dishes, full of incense, weighing 10 shekels apiece according to the shekel of the sanctuary, all the gold of the dishes being 120 shekels;
NUM|7|87|all the cattle for the burnt offering twelve bulls, twelve rams, twelve male lambs a year old, with their grain offering; and twelve male goats for a sin offering;
NUM|7|88|and all the cattle for the sacrifice of peace offerings twenty-four bulls, the rams sixty, the male goats sixty, the male lambs a year old sixty. This was the dedication offering for the altar after it was anointed.
NUM|7|89|And when Moses went into the tent of meeting to speak with the LORD, he heard the voice speaking to him from above the mercy seat that was on the ark of the testimony, from between the two cherubim; and it spoke to him.
NUM|8|1|Now the LORD spoke to Moses, saying,
NUM|8|2|"Speak to Aaron and say to him, When you set up the lamps, the seven lamps shall give light in front of the lampstand."
NUM|8|3|And Aaron did so: he set up its lamps in front of the lampstand, as the LORD commanded Moses.
NUM|8|4|And this was the workmanship of the lampstand, hammered work of gold. From its base to its flowers, it was hammered work; according to the pattern that the LORD had shown Moses, so he made the lampstand.
NUM|8|5|And the LORD spoke to Moses, saying,
NUM|8|6|"Take the Levites from among the people of Israel and cleanse them.
NUM|8|7|Thus you shall do to them to cleanse them: sprinkle the water of purification upon them, and let them go with a razor over all their body, and wash their clothes and cleanse themselves.
NUM|8|8|Then let them take a bull from the herd and its grain offering of fine flour mixed with oil, and you shall take another bull from the herd for a sin offering.
NUM|8|9|And you shall bring the Levites before the tent of meeting and assemble the whole congregation of the people of Israel.
NUM|8|10|When you bring the Levites before the LORD, the people of Israel shall lay their hands on the Levites,
NUM|8|11|and Aaron shall offer the Levites before the LORD as a wave offering from the people of Israel, that they may do the service of the LORD.
NUM|8|12|Then the Levites shall lay their hands on the heads of the bulls, and you shall offer the one for a sin offering and the other for a burnt offering to the LORD to make atonement for the Levites.
NUM|8|13|And you shall set the Levites before Aaron and his sons, and shall offer them as a wave offering to the LORD.
NUM|8|14|"Thus you shall separate the Levites from among the people of Israel, and the Levites shall be mine.
NUM|8|15|And after that the Levites shall go in to serve at the tent of meeting, when you have cleansed them and offered them as a wave offering.
NUM|8|16|For they are wholly given to me from among the people of Israel. Instead of all who open the womb, the firstborn of all the people of Israel, I have taken them for myself.
NUM|8|17|For all the firstborn among the people of Israel are mine, both of man and of beast. On the day that I struck down all the firstborn in the land of Egypt I consecrated them for myself,
NUM|8|18|and I have taken the Levites instead of all the firstborn among the people of Israel.
NUM|8|19|And I have given the Levites as a gift to Aaron and his sons from among the people of Israel, to do the service for the people of Israel at the tent of meeting and to make atonement for the people of Israel, that there may be no plague among the people of Israel when the people of Israel come near the sanctuary."
NUM|8|20|Thus did Moses and Aaron and all the congregation of the people of Israel to the Levites. According to all that the LORD commanded Moses concerning the Levites, the people of Israel did to them.
NUM|8|21|And the Levites purified themselves from sin and washed their clothes, and Aaron offered them as a wave offering before the LORD, and Aaron made atonement for them to cleanse them.
NUM|8|22|And after that the Levites went in to do their service in the tent of meeting before Aaron and his sons; as the LORD had commanded Moses concerning the Levites, so they did to them.
NUM|8|23|And the LORD spoke to Moses, saying,
NUM|8|24|"This applies to the Levites: from twenty-five years old and upward they shall come to do duty in the service of the tent of meeting.
NUM|8|25|And from the age of fifty years they shall withdraw from the duty of the service and serve no more.
NUM|8|26|They minister to their brothers in the tent of meeting by keeping guard, but they shall do no service. Thus shall you do to the Levites in assigning their duties."
NUM|9|1|And the LORD spoke to Moses in the wilderness of Sinai, in the first month of the second year after they had come out of the land of Egypt, saying,
NUM|9|2|"Let the people of Israel keep the Passover at its appointed time.
NUM|9|3|On the fourteenth day of this month, at twilight, you shall keep it at its appointed time; according to all its statutes and all its rules you shall keep it."
NUM|9|4|So Moses told the people of Israel that they should keep the Passover.
NUM|9|5|And they kept the Passover in the first month, on the fourteenth day of the month, at twilight, in the wilderness of Sinai; according to all that the LORD commanded Moses, so the people of Israel did.
NUM|9|6|And there were certain men who were unclean through touching a dead body, so that they could not keep the Passover on that day, and they came before Moses and Aaron on that day.
NUM|9|7|And those men said to him, "We are unclean through touching a dead body. Why are we kept from bringing the LORD's offering at its appointed time among the people of Israel?"
NUM|9|8|And Moses said to them, "Wait, that I may hear what the LORD will command concerning you."
NUM|9|9|The LORD spoke to Moses, saying,
NUM|9|10|"Speak to the people of Israel, saying, If any one of you or of your descendants is unclean through touching a dead body, or is on a long journey, he shall still keep the Passover to the LORD.
NUM|9|11|In the second month on the fourteenth day at twilight they shall keep it. They shall eat it with unleavened bread and bitter herbs.
NUM|9|12|They shall leave none of it until the morning, nor break any of its bones; according to all the statute for the Passover they shall keep it.
NUM|9|13|But if anyone who is clean and is not on a journey fails to keep the Passover, that person shall be cut off from his people because he did not bring the LORD's offering at its appointed time; that man shall bear his sin.
NUM|9|14|And if a stranger sojourns among you and would keep the Passover to the LORD, according to the statute of the Passover and according to its rule, so shall he do. You shall have one statute, both for the sojourner and for the native."
NUM|9|15|On the day that the tabernacle was set up, the cloud covered the tabernacle, the tent of the testimony. And at evening it was over the tabernacle like the appearance of fire until morning.
NUM|9|16|So it was always: the cloud covered it by day and the appearance of fire by night.
NUM|9|17|And whenever the cloud lifted from over the tent, after that the people of Israel set out, and in the place where the cloud settled down, there the people of Israel camped.
NUM|9|18|At the command of the LORD the people of Israel set out, and at the command of the LORD they camped. As long as the cloud rested over the tabernacle, they remained in camp.
NUM|9|19|Even when the cloud continued over the tabernacle many days, the people of Israel kept the charge of the LORD and did not set out.
NUM|9|20|Sometimes the cloud was a few days over the tabernacle, and according to the command of the LORD they remained in camp; then according to the command of the LORD they set out.
NUM|9|21|And sometimes the cloud remained from evening until morning. And when the cloud lifted in the morning, they set out, or if it continued for a day and a night, when the cloud lifted they set out.
NUM|9|22|Whether it was two days, or a month, or a longer time, that the cloud continued over the tabernacle, abiding there, the people of Israel remained in camp and did not set out, but when it lifted they set out.
NUM|9|23|At the command of the LORD they camped, and at the command of the LORD they set out. They kept the charge of the LORD, at the command of the LORD by Moses.
NUM|10|1|The LORD spoke to Moses, saying,
NUM|10|2|"Make two silver trumpets. Of hammered work you shall make them, and you shall use them for summoning the congregation and for breaking camp.
NUM|10|3|And when both are blown, all the congregation shall gather themselves to you at the entrance of the tent of meeting.
NUM|10|4|But if they blow only one, then the chiefs, the heads of the tribes of Israel, shall gather themselves to you.
NUM|10|5|When you blow an alarm, the camps that are on the east side shall set out.
NUM|10|6|And when you blow an alarm the second time, the camps that are on the south side shall set out. An alarm is to be blown whenever they are to set out.
NUM|10|7|But when the assembly is to be gathered together, you shall blow a long blast, but you shall not sound an alarm.
NUM|10|8|And the sons of Aaron, the priests, shall blow the trumpets. The trumpets shall be to you for a perpetual statute throughout your generations.
NUM|10|9|And when you go to war in your land against the adversary who oppresses you, then you shall sound an alarm with the trumpets, that you may be remembered before the LORD your God, and you shall be saved from your enemies.
NUM|10|10|On the day of your gladness also, and at your appointed feasts and at the beginnings of your months, you shall blow the trumpets over your burnt offerings and over the sacrifices of your peace offerings. They shall be a reminder of you before your God: I am the LORD your God."
NUM|10|11|In the second year, in the second month, on the twentieth day of the month, the cloud lifted from over the tabernacle of the testimony,
NUM|10|12|and the people of Israel set out by stages from the wilderness of Sinai. And the cloud settled down in the wilderness of Paran.
NUM|10|13|They set out for the first time at the command of the LORD by Moses.
NUM|10|14|The standard of the camp of the people of Judah set out first by their companies, and over their company was Nahshon the son of Amminadab.
NUM|10|15|And over the company of the tribe of the people of Issachar was Nethanel the son of Zuar.
NUM|10|16|And over the company of the tribe of the people of Zebulun was Eliab the son of Helon.
NUM|10|17|And when the tabernacle was taken down, the sons of Gershon and the sons of Merari, who carried the tabernacle, set out.
NUM|10|18|And the standard of the camp of Reuben set out by their companies, and over their company was Elizur the son of Shedeur.
NUM|10|19|And over the company of the tribe of the people of Simeon was Shelumiel the son of Zurishaddai.
NUM|10|20|And over the company of the tribe of the people of Gad was Eliasaph the son of Deuel.
NUM|10|21|Then the Kohathites set out, carrying the holy things, and the tabernacle was set up before their arrival.
NUM|10|22|And the standard of the camp of the people of Ephraim set out by their companies, and over their company was Elishama the son of Ammihud.
NUM|10|23|And over the company of the tribe of the people of Manasseh was Gamaliel the son of Pedahzur.
NUM|10|24|And over the company of the tribe of the people of Benjamin was Abidan the son of Gideoni.
NUM|10|25|Then the standard of the camp of the people of Dan, acting as the rear guard of all the camps, set out by their companies, and over their company was Ahiezer the son of Ammishaddai.
NUM|10|26|And over the company of the tribe of the people of Asher was Pagiel the son of Ochran.
NUM|10|27|And over the company of the tribe of the people of Naphtali was Ahira the son of Enan.
NUM|10|28|This was the order of march of the people of Israel by their companies, when they set out.
NUM|10|29|And Moses said to Hobab the son of Reuel the Midianite, Moses' father-in-law, "We are setting out for the place of which the LORD said, 'I will give it to you.' Come with us, and we will do good to you, for the LORD has promised good to Israel."
NUM|10|30|But he said to him, "I will not go. I will depart to my own land and to my kindred."
NUM|10|31|And he said, "Please do not leave us, for you know where we should camp in the wilderness, and you will serve as eyes for us.
NUM|10|32|And if you do go with us, whatever good the LORD will do to us, the same will we do to you."
NUM|10|33|So they set out from the mount of the LORD three days' journey. And the ark of the covenant of the LORD went before them three days' journey, to seek out a resting place for them.
NUM|10|34|And the cloud of the LORD was over them by day, whenever they set out from the camp.
NUM|10|35|And whenever the ark set out, Moses said, "Arise, O LORD, and let your enemies be scattered, and let those who hate you flee before you."
NUM|10|36|And when it rested, he said, "Return, O LORD, to the ten thousand thousands of Israel."
NUM|11|1|And the people complained in the hearing of the LORD about their misfortunes, and when the LORD heard it, his anger was kindled, and the fire of the LORD burned among them and consumed some outlying parts of the camp.
NUM|11|2|Then the people cried out to Moses, and Moses prayed to the LORD, and the fire died down.
NUM|11|3|So the name of that place was called Taberah, because the fire of the LORD burned among them.
NUM|11|4|Now the rabble that was among them had a strong craving. And the people of Israel also wept again and said, "Oh that we had meat to eat!
NUM|11|5|We remember the fish we ate in Egypt that cost nothing, the cucumbers, the melons, the leeks, the onions, and the garlic.
NUM|11|6|But now our strength is dried up, and there is nothing at all but this manna to look at."
NUM|11|7|Now the manna was like coriander seed, and its appearance like that of bdellium.
NUM|11|8|The people went about and gathered it and ground it in hand-mills or beat it in mortars and boiled it in pots and made cakes of it. And the taste of it was like the taste of cakes baked with oil.
NUM|11|9|When the dew fell upon the camp in the night, the manna fell with it.
NUM|11|10|Moses heard the people weeping throughout their clans, everyone at the door of his tent. And the anger of the LORD blazed hotly, and Moses was displeased.
NUM|11|11|Moses said to the LORD, "Why have you dealt ill with your servant? And why have I not found favor in your sight, that you lay the burden of all this people on me?
NUM|11|12|Did I conceive all this people? Did I give them birth, that you should say to me, 'Carry them in your bosom, as a nurse carries a nursing child,' to the land that you swore to give their fathers?
NUM|11|13|Where am I to get meat to give to all this people? For they weep before me and say, 'Give us meat, that we may eat.'
NUM|11|14|I am not able to carry all this people alone; the burden is too heavy for me.
NUM|11|15|If you will treat me like this, kill me at once, if I find favor in your sight, that I may not see my wretchedness."
NUM|11|16|Then the LORD said to Moses, "Gather for me seventy men of the elders of Israel, whom you know to be the elders of the people and officers over them, and bring them to the tent of meeting, and let them take their stand there with you.
NUM|11|17|And I will come down and talk with you there. And I will take some of the Spirit that is on you and put it on them, and they shall bear the burden of the people with you, so that you may not bear it yourself alone.
NUM|11|18|And say to the people, 'Consecrate yourselves for tomorrow, and you shall eat meat, for you have wept in the hearing of the LORD, saying, "Who will give us meat to eat? For it was better for us in Egypt." Therefore the LORD will give you meat, and you shall eat.
NUM|11|19|You shall not eat just one day, or two days, or five days, or ten days, or twenty days,
NUM|11|20|but a whole month, until it comes out at your nostrils and becomes loathsome to you, because you have rejected the LORD who is among you and have wept before him, saying, "Why did we come out of Egypt?"'"
NUM|11|21|But Moses said, "The people among whom I am number six hundred thousand on foot, and you have said, 'I will give them meat, that they may eat a whole month!'
NUM|11|22|Shall flocks and herds be slaughtered for them, and be enough for them? Or shall all the fish of the sea be gathered together for them, and be enough for them?"
NUM|11|23|And the LORD said to Moses, "Is the LORD's hand shortened? Now you shall see whether my word will come true for you or not."
NUM|11|24|So Moses went out and told the people the words of the LORD. And he gathered seventy men of the elders of the people and placed them around the tent.
NUM|11|25|Then the LORD came down in the cloud and spoke to him, and took some of the Spirit that was on him and put it on the seventy elders. And as soon as the Spirit rested on them, they prophesied. But they did not continue doing it.
NUM|11|26|Now two men remained in the camp, one named Eldad, and the other named Medad, and the Spirit rested on them. They were among those registered, but they had not gone out to the tent, and so they prophesied in the camp.
NUM|11|27|And a young man ran and told Moses, "Eldad and Medad are prophesying in the camp."
NUM|11|28|And Joshua the son of Nun, the assistant of Moses from his youth, said, "My lord Moses, stop them."
NUM|11|29|But Moses said to him, "Are you jealous for my sake? Would that all the LORD's people were prophets, that the LORD would put his Spirit on them!"
NUM|11|30|And Moses and the elders of Israel returned to the camp.
NUM|11|31|Then a wind from the LORD sprang up, and it brought quail from the sea and let them fall beside the camp, about a day's journey on this side and a day's journey on the other side, around the camp, and about two cubits above the ground.
NUM|11|32|And the people rose all that day and all night and all the next day, and gathered the quail. Those who gathered least gathered ten homers. And they spread them out for themselves all around the camp.
NUM|11|33|While the meat was yet between their teeth, before it was consumed, the anger of the LORD was kindled against the people, and the LORD struck down the people with a very great plague.
NUM|11|34|Therefore the name of that place was called Kibroth-hattaavah, because there they buried the people who had the craving.
NUM|11|35|From Kibroth-hattaavah the people journeyed to Hazeroth, and they remained at Hazeroth.
NUM|12|1|Miriam and Aaron spoke against Moses because of the Cushite woman whom he had married, for he had married a Cushite woman.
NUM|12|2|And they said, "Has the LORD indeed spoken only through Moses? Has he not spoken through us also?" And the LORD heard it.
NUM|12|3|Now the man Moses was very meek, more than all people who were on the face of the earth.
NUM|12|4|And suddenly the LORD said to Moses and to Aaron and Miriam, "Come out, you three, to the tent of meeting." And the three of them came out.
NUM|12|5|And the LORD came down in a pillar of cloud and stood at the entrance of the tent and called Aaron and Miriam, and they both came forward.
NUM|12|6|And he said, "Hear my words: If there is a prophet among you, I the LORD make myself known to him in a vision; I speak with him in a dream.
NUM|12|7|Not so with my servant Moses. He is faithful in all my house.
NUM|12|8|With him I speak mouth to mouth, clearly, and not in riddles, and he beholds the form of the LORD. Why then were you not afraid to speak against my servant Moses?"
NUM|12|9|And the anger of the LORD was kindled against them, and he departed.
NUM|12|10|When the cloud removed from over the tent, behold, Miriam was leprous, like snow. And Aaron turned toward Miriam, and behold, she was leprous.
NUM|12|11|And Aaron said to Moses, "Oh, my lord, do not punish us because we have done foolishly and have sinned.
NUM|12|12|Let her not be as one dead, whose flesh is half eaten away when he comes out of his mother's womb."
NUM|12|13|And Moses cried to the LORD, "O God, please heal her- please."
NUM|12|14|But the LORD said to Moses, "If her father had but spit in her face, should she not be shamed seven days? Let her be shut outside the camp seven days, and after that she may be brought in again."
NUM|12|15|So Miriam was shut outside the camp seven days, and the people did not set out on the march till Miriam was brought in again.
NUM|12|16|After that the people set out from Hazeroth, and camped in the wilderness of Paran.
NUM|13|1|The LORD spoke to Moses, saying,
NUM|13|2|"Send men to spy out the land of Canaan, which I am giving to the people of Israel. From each tribe of their fathers you shall send a man, every one a chief among them."
NUM|13|3|So Moses sent them from the wilderness of Paran, according to the command of the LORD, all of them men who were heads of the people of Israel.
NUM|13|4|And these were their names: From the tribe of Reuben, Shammua the son of Zaccur;
NUM|13|5|from the tribe of Simeon, Shaphat the son of Hori;
NUM|13|6|from the tribe of Judah, Caleb the son of Jephunneh;
NUM|13|7|from the tribe of Issachar, Igal the son of Joseph;
NUM|13|8|from the tribe of Ephraim, Hoshea the son of Nun;
NUM|13|9|from the tribe of Benjamin, Palti the son of Raphu;
NUM|13|10|from the tribe of Zebulun, Gaddiel the son of Sodi;
NUM|13|11|from the tribe of Joseph (that is, from the tribe of Manasseh), Gaddi the son of Susi;
NUM|13|12|from the tribe of Dan, Ammiel the son of Gemalli;
NUM|13|13|from the tribe of Asher, Sethur the son of Michael;
NUM|13|14|from the tribe of Naphtali, Nahbi the son of Vophsi;
NUM|13|15|from the tribe of Gad, Geuel the son of Machi.
NUM|13|16|These were the names of the men whom Moses sent to spy out the land. And Moses called Hoshea the son of Nun Joshua.
NUM|13|17|Moses sent them to spy out the land of Canaan and said to them, "Go up into the Negeb and go up into the hill country,
NUM|13|18|and see what the land is, and whether the people who dwell in it are strong or weak, whether they are few or many,
NUM|13|19|and whether the land that they dwell in is good or bad, and whether the cities that they dwell in are camps or strongholds,
NUM|13|20|and whether the land is rich or poor, and whether there are trees in it or not. Be of good courage and bring some of the fruit of the land." Now the time was the season of the first ripe grapes.
NUM|13|21|So they went up and spied out the land from the wilderness of Zin to Rehob, near Lebo-hamath.
NUM|13|22|They went up into the Negeb and came to Hebron. Ahiman, Sheshai, and Talmai, the descendants of Anak, were there. (Hebron was built seven years before Zoan in Egypt.)
NUM|13|23|And they came to the Valley of Eshcol and cut down from there a branch with a single cluster of grapes, and they carried it on a pole between two of them; they also brought some pomegranates and figs.
NUM|13|24|That place was called the Valley of Eshcol, because of the cluster that the people of Israel cut down from there.
NUM|13|25|At the end of forty days they returned from spying out the land.
NUM|13|26|And they came to Moses and Aaron and to all the congregation of the people of Israel in the wilderness of Paran, at Kadesh. They brought back word to them and to all the congregation, and showed them the fruit of the land.
NUM|13|27|And they told him, "We came to the land to which you sent us. It flows with milk and honey, and this is its fruit.
NUM|13|28|However, the people who dwell in the land are strong, and the cities are fortified and very large. And besides, we saw the descendants of Anak there.
NUM|13|29|The Amalekites dwell in the land of the Negeb. The Hittites, the Jebusites, and the Amorites dwell in the hill country. And the Canaanites dwell by the sea, and along the Jordan."
NUM|13|30|But Caleb quieted the people before Moses and said, "Let us go up at once and occupy it, for we are well able to overcome it."
NUM|13|31|Then the men who had gone up with him said, "We are not able to go up against the people, for they are stronger than we are."
NUM|13|32|So they brought to the people of Israel a bad report of the land that they had spied out, saying, "The land, through which we have gone to spy it out, is a land that devours its inhabitants, and all the people that we saw in it are of great height.
NUM|13|33|And there we saw the Nephilim (the sons of Anak, who come from the Nephilim), and we seemed to ourselves like grasshoppers, and so we seemed to them."
NUM|14|1|Then all the congregation raised a loud cry, and the people wept that night.
NUM|14|2|And all the people of Israel grumbled against Moses and Aaron. The whole congregation said to them, "Would that we had died in the land of Egypt! Or would that we had died in this wilderness!
NUM|14|3|Why is the LORD bringing us into this land, to fall by the sword? Our wives and our little ones will become a prey. Would it not be better for us to go back to Egypt?"
NUM|14|4|And they said to one another, "Let us choose a leader and go back to Egypt."
NUM|14|5|Then Moses and Aaron fell on their faces before all the assembly of the congregation of the people of Israel.
NUM|14|6|And Joshua the son of Nun and Caleb the son of Jephunneh, who were among those who had spied out the land, tore their clothes
NUM|14|7|and said to all the congregation of the people of Israel, "The land, which we passed through to spy it out, is an exceedingly good land.
NUM|14|8|If the LORD delights in us, he will bring us into this land and give it to us, a land that flows with milk and honey.
NUM|14|9|Only do not rebel against the LORD. And do not fear the people of the land, for they are bread for us. Their protection is removed from them, and the LORD is with us; do not fear them."
NUM|14|10|Then all the congregation said to stone them with stones. But the glory of the LORD appeared at the tent of meeting to all the people of Israel.
NUM|14|11|And the LORD said to Moses, "How long will this people despise me? And how long will they not believe in me, in spite of all the signs that I have done among them?
NUM|14|12|I will strike them with the pestilence and disinherit them, and I will make of you a nation greater and mightier than they."
NUM|14|13|But Moses said to the LORD, "Then the Egyptians will hear of it, for you brought up this people in your might from among them,
NUM|14|14|and they will tell the inhabitants of this land. They have heard that you, O LORD, are in the midst of this people. For you, O LORD, are seen face to face, and your cloud stands over them and you go before them, in a pillar of cloud by day and in a pillar of fire by night.
NUM|14|15|Now if you kill this people as one man, then the nations who have heard your fame will say,
NUM|14|16|'It is because the LORD was not able to bring this people into the land that he swore to give to them that he has killed them in the wilderness.'
NUM|14|17|And now, please let the power of the Lord be great as you have promised, saying,
NUM|14|18|'The LORD is slow to anger and abounding in steadfast love, forgiving iniquity and transgression, but he will by no means clear the guilty, visiting the iniquity of the fathers on the children, to the third and the fourth generation.'
NUM|14|19|Please pardon the iniquity of this people, according to the greatness of your steadfast love, just as you have forgiven this people, from Egypt until now."
NUM|14|20|Then the LORD said, "I have pardoned, according to your word.
NUM|14|21|But truly, as I live, and as all the earth shall be filled with the glory of the LORD,
NUM|14|22|none of the men who have seen my glory and my signs that I did in Egypt and in the wilderness, and yet have put me to the test these ten times and have not obeyed my voice,
NUM|14|23|shall see the land that I swore to give to their fathers. And none of those who despised me shall see it.
NUM|14|24|But my servant Caleb, because he has a different spirit and has followed me fully, I will bring into the land into which he went, and his descendants shall possess it.
NUM|14|25|Now, since the Amalekites and the Canaanites dwell in the valleys, turn tomorrow and set out for the wilderness by the way to the Red Sea."
NUM|14|26|And the LORD spoke to Moses and to Aaron, saying,
NUM|14|27|"How long shall this wicked congregation grumble against me? I have heard the grumblings of the people of Israel, which they grumble against me.
NUM|14|28|Say to them, 'As I live, declares the LORD, what you have said in my hearing I will do to you:
NUM|14|29|your dead bodies shall fall in this wilderness, and of all your number, listed in the census from twenty years old and upward, who have grumbled against me,
NUM|14|30|not one shall come into the land where I swore that I would make you dwell, except Caleb the son of Jephunneh and Joshua the son of Nun.
NUM|14|31|But your little ones, who you said would become a prey, I will bring in, and they shall know the land that you have rejected.
NUM|14|32|But as for you, your dead bodies shall fall in this wilderness.
NUM|14|33|And your children shall be shepherds in the wilderness forty years and shall suffer for your faithlessness, until the last of your dead bodies lies in the wilderness.
NUM|14|34|According to the number of the days in which you spied out the land, forty days, a year for each day, you shall bear your iniquity forty years, and you shall know my displeasure.'
NUM|14|35|I, the LORD, have spoken. Surely this will I do to all this wicked congregation who are gathered together against me: in this wilderness they shall come to a full end, and there they shall die."
NUM|14|36|And the men whom Moses sent to spy out the land, who returned and made all the congregation grumble against him by bringing up a bad report about the land-
NUM|14|37|the men who brought up a bad report of the land- died by plague before the LORD.
NUM|14|38|Of those men who went to spy out the land, only Joshua the son of Nun and Caleb the son of Jephunneh remained alive.
NUM|14|39|When Moses told these words to all the people of Israel, the people mourned greatly.
NUM|14|40|And they rose early in the morning and went up to the heights of the hill country, saying, "Here we are. We will go up to the place that the LORD has promised, for we have sinned."
NUM|14|41|But Moses said, "Why now are you transgressing the command of the LORD, when that will not succeed?
NUM|14|42|Do not go up, for the Lord is not among you, lest you be struck down before your enemies.
NUM|14|43|For there the Amalekites and the Canaanites are facing you, and you shall fall by the sword. Because you have turned back from following the LORD, the LORD will not be with you."
NUM|14|44|But they presumed to go up to the heights of the hill country, although neither the ark of the covenant of the LORD nor Moses departed out of the camp.
NUM|14|45|Then the Amalekites and the Canaanites who lived in that hill country came down and defeated them and pursued them, even to Hormah.
NUM|15|1|The LORD spoke to Moses, saying,
NUM|15|2|"Speak to the people of Israel and say to them, When you come into the land you are to inhabit, which I am giving you,
NUM|15|3|and you offer to the LORD from the herd or from the flock a food offering or a burnt offering or a sacrifice, to fulfill a vow or as a freewill offering or at your appointed feasts, to make a pleasing aroma to the LORD,
NUM|15|4|then he who brings his offering shall offer to the LORD a grain offering of a tenth of an ephah of fine flour, mixed with a quarter of a hin of oil;
NUM|15|5|and you shall offer with the burnt offering, or for the sacrifice, a quarter of a hin of wine for the drink offering for each lamb.
NUM|15|6|Or for a ram, you shall offer for a grain offering two tenths of an ephah of fine flour mixed with a third of a hin of oil.
NUM|15|7|And for the drink offering you shall offer a third of a hin of wine, a pleasing aroma to the LORD.
NUM|15|8|And when you offer a bull as a burnt offering or sacrifice, to fulfill a vow or for peace offerings to the LORD,
NUM|15|9|then one shall offer with the bull a grain offering of three tenths of an ephah of fine flour, mixed with half a hin of oil.
NUM|15|10|And you shall offer for the drink offering half a hin of wine, as a food offering, a pleasing aroma to the LORD.
NUM|15|11|"Thus it shall be done for each bull or ram, or for each lamb or young goat.
NUM|15|12|As many as you offer, so shall you do with each one, as many as there are.
NUM|15|13|Every native Israelite shall do these things in this way, in offering a food offering, with a pleasing aroma to the LORD.
NUM|15|14|And if a stranger is sojourning with you, or anyone is living permanently among you, and he wishes to offer a food offering, with a pleasing aroma to the LORD, he shall do as you do.
NUM|15|15|For the assembly, there shall be one statute for you and for the stranger who sojourns with you, a statute forever throughout your generations. You and the sojourner shall be alike before the LORD.
NUM|15|16|One law and one rule shall be for you and for the stranger who sojourns with you."
NUM|15|17|The LORD spoke to Moses, saying,
NUM|15|18|"Speak to the people of Israel and say to them, When you come into the land to which I bring you
NUM|15|19|and when you eat of the bread of the land, you shall present a contribution to the LORD.
NUM|15|20|Of the first of your dough you shall present a loaf as a contribution; like a contribution from the threshing floor, so shall you present it.
NUM|15|21|Some of the first of your dough you shall give to the LORD as a contribution throughout your generations.
NUM|15|22|"But if you sin unintentionally, and do not observe all these commandments that the LORD has spoken to Moses,
NUM|15|23|all that the LORD has commanded you by Moses, from the day that the LORD gave commandment, and onward throughout your generations,
NUM|15|24|then if it was done unintentionally without the knowledge of the congregation, all the congregation shall offer one bull from the herd for a burnt offering, a pleasing aroma to the LORD, with its grain offering and its drink offering, according to the rule, and one male goat for a sin offering.
NUM|15|25|And the priest shall make atonement for all the congregation of the people of Israel, and they shall be forgiven, because it was a mistake, and they have brought their offering, a food offering to the LORD, and their sin offering before the LORD for their mistake.
NUM|15|26|And all the congregation of the people of Israel shall be forgiven, and the stranger who sojourns among them, because the whole population was involved in the mistake.
NUM|15|27|"If one person sins unintentionally, he shall offer a female goat a year old for a sin offering.
NUM|15|28|And the priest shall make atonement before the LORD for the person who makes a mistake, when he sins unintentionally, to make atonement for him, and he shall be forgiven.
NUM|15|29|You shall have one law for him who does anything unintentionally, for him who is native among the people of Israel and for the stranger who sojourns among them.
NUM|15|30|But the person who does anything with a high hand, whether he is native or a sojourner, reviles the LORD, and that person shall be cut off from among his people.
NUM|15|31|Because he has despised the word of the LORD and has broken his commandment, that person shall be utterly cut off; his iniquity shall be on him."
NUM|15|32|While the people of Israel were in the wilderness, they found a man gathering sticks on the Sabbath day.
NUM|15|33|And those who found him gathering sticks brought him to Moses and Aaron and to all the congregation.
NUM|15|34|They put him in custody, because it had not been made clear what should be done to him.
NUM|15|35|And the LORD said to Moses, "The man shall be put to death; all the congregation shall stone him with stones outside the camp."
NUM|15|36|And all the congregation brought him outside the camp and stoned him to death with stones, as the LORD commanded Moses.
NUM|15|37|The LORD said to Moses,
NUM|15|38|"Speak to the people of Israel, and tell them to make tassels on the corners of their garments throughout their generations, and to put a cord of blue on the tassel of each corner.
NUM|15|39|And it shall be a tassel for you to look at and remember all the commandments of the LORD, to do them, not to follow after your own heart and your own eyes, which you are inclined to whore after.
NUM|15|40|So you shall remember and do all my commandments, and be holy to your God.
NUM|15|41|I am the LORD your God, who brought you out of the land of Egypt to be your God: I am the LORD your God."
NUM|16|1|Now Korah the son of Izhar, son of Kohath, son of Levi, and Dathan and Abiram the sons of Eliab, and On the son of Peleth, sons of Reuben, took men.
NUM|16|2|And they rose up before Moses, with a number of the people of Israel, 250 chiefs of the congregation, chosen from the assembly, well-known men.
NUM|16|3|They assembled themselves together against Moses and against Aaron and said to them, "You have gone too far! For all in the congregation are holy, every one of them, and the LORD is among them. Why then do you exalt yourselves above the assembly of the LORD?"
NUM|16|4|When Moses heard it, he fell on his face,
NUM|16|5|and he said to Korah and all his company, "In the morning the LORD will show who is his, and who is holy, and will bring him near to him. The one whom he chooses he will bring near to him.
NUM|16|6|Do this: take censers, Korah and all his company;
NUM|16|7|put fire in them and put incense on them before the LORD tomorrow, and the man whom the LORD chooses shall be the holy one. You have gone too far, sons of Levi!"
NUM|16|8|And Moses said to Korah, "Hear now, you sons of Levi:
NUM|16|9|is it too small a thing for you that the God of Israel has separated you from the congregation of Israel, to bring you near to himself, to do service in the tabernacle of the LORD and to stand before the congregation to minister to them,
NUM|16|10|and that he has brought you near him, and all your brothers the sons of Levi with you? And would you seek the priesthood also?
NUM|16|11|Therefore it is against the LORD that you and all your company have gathered together. What is Aaron that you grumble against him?"
NUM|16|12|And Moses sent to call Dathan and Abiram the sons of Eliab, and they said, "We will not come up.
NUM|16|13|Is it a small thing that you have brought us up out of a land flowing with milk and honey, to kill us in the wilderness, that you must also make yourself a prince over us?
NUM|16|14|Moreover, you have not brought us into a land flowing with milk and honey, nor given us inheritance of fields and vineyards. Will you put out the eyes of these men? We will not come up."
NUM|16|15|And Moses was very angry and said to the LORD, "Do not respect their offering. I have not taken one donkey from them, and I have not harmed one of them."
NUM|16|16|And Moses said to Korah, "Be present, you and all your company, before the LORD, you and they, and Aaron, tomorrow.
NUM|16|17|And let every one of you take his censer and put incense on it, and every one of you bring before the LORD his censer, 250 censers; you also, and Aaron, each his censer."
NUM|16|18|So every man took his censer and put fire in them and laid incense on them and stood at the entrance of the tent of meeting with Moses and Aaron.
NUM|16|19|Then Korah assembled all the congregation against them at the entrance of the tent of meeting. And the glory of the LORD appeared to all the congregation.
NUM|16|20|And the LORD spoke to Moses and to Aaron, saying,
NUM|16|21|"Separate yourselves from among this congregation, that I may consume them in a moment."
NUM|16|22|And they fell on their faces and said, "O God, the God of the spirits of all flesh, shall one man sin, and will you be angry with all the congregation?"
NUM|16|23|And the LORD spoke to Moses, saying,
NUM|16|24|"Say to the congregation, Get away from the dwelling of Korah, Dathan, and Abiram."
NUM|16|25|Then Moses rose and went to Dathan and Abiram, and the elders of Israel followed him.
NUM|16|26|And he spoke to the congregation, saying, "Depart, please, from the tents of these wicked men, and touch nothing of theirs, lest you be swept away with all their sins."
NUM|16|27|So they got away from the dwelling of Korah, Dathan, and Abiram. And Dathan and Abiram came out and stood at the door of their tents, together with their wives, their sons, and their little ones.
NUM|16|28|And Moses said, "Hereby you shall know that the LORD has sent me to do all these works, and that it has not been of my own accord.
NUM|16|29|If these men die as all men die, or if they are visited by the fate of all mankind, then the LORD has not sent me.
NUM|16|30|But if the LORD creates something new, and the ground opens its mouth and swallows them up with all that belongs to them, and they go down alive into Sheol, then you shall know that these men have despised the LORD."
NUM|16|31|And as soon as he had finished speaking all these words, the ground under them split apart.
NUM|16|32|And the earth opened its mouth and swallowed them up, with their households and all the people who belonged to Korah and all their goods.
NUM|16|33|So they and all that belonged to them went down alive into Sheol, and the earth closed over them, and they perished from the midst of the assembly.
NUM|16|34|And all Israel who were around them fled at their cry, for they said, "Lest the earth swallow us up!"
NUM|16|35|And fire came out from the LORD and consumed the 250 men offering the incense.
NUM|16|36|Then the LORD spoke to Moses, saying,
NUM|16|37|"Tell Eleazar the son of Aaron the priest to take up the censers out of the blaze. Then scatter the fire far and wide, for they have become holy.
NUM|16|38|As for the censers of these men who have sinned at the cost of their lives, let them be made into hammered plates as a covering for the altar, for they offered them before the LORD, and they became holy. Thus they shall be a sign to the people of Israel."
NUM|16|39|So Eleazar the priest took the bronze censers, which those who were burned had offered, and they were hammered out as a covering for the altar,
NUM|16|40|to be a reminder to the people of Israel, so that no outsider, who is not of the descendants of Aaron, should draw near to burn incense before the LORD, lest he become like Korah and his company- as the LORD said to him through Moses.
NUM|16|41|But on the next day all the congregation of the people of Israel grumbled against Moses and against Aaron, saying, "You have killed the people of the LORD."
NUM|16|42|And when the congregation had assembled against Moses and against Aaron, they turned toward the tent of meeting. And behold, the cloud covered it, and the glory of the LORD appeared.
NUM|16|43|And Moses and Aaron came to the front of the tent of meeting,
NUM|16|44|and the LORD spoke to Moses, saying,
NUM|16|45|"Get away from the midst of this congregation, that I may consume them in a moment." And they fell on their faces.
NUM|16|46|And Moses said to Aaron, "Take your censer, and put fire on it from off the altar and lay incense on it and carry it quickly to the congregation and make atonement for them, for wrath has gone out from the LORD; the plague has begun."
NUM|16|47|So Aaron took it as Moses said and ran into the midst of the assembly. And behold, the plague had already begun among the people. And he put on the incense and made atonement for the people.
NUM|16|48|And he stood between the dead and the living, and the plague was stopped.
NUM|16|49|Now those who died in the plague were 14,700, besides those who died in the affair of Korah.
NUM|16|50|And Aaron returned to Moses at the entrance of the tent of meeting, when the plague was stopped.
NUM|17|1|The LORD spoke to Moses, saying,
NUM|17|2|"Speak to the people of Israel, and get from them staffs, one for each fathers' house, from all their chiefs according to their fathers' houses, twelve staffs. Write each man's name on his staff,
NUM|17|3|and write Aaron's name on the staff of Levi. For there shall be one staff for the head of each fathers' house.
NUM|17|4|Then you shall deposit them in the tent of meeting before the testimony, where I meet with you.
NUM|17|5|And the staff of the man whom I choose shall sprout. Thus I will make to cease from me the grumblings of the people of Israel, which they grumble against you."
NUM|17|6|Moses spoke to the people of Israel. And all their chiefs gave him staffs, one for each chief, according to their fathers' houses, twelve staffs. And the staff of Aaron was among their staffs.
NUM|17|7|And Moses deposited the staffs before the LORD in the tent of the testimony.
NUM|17|8|On the next day Moses went into the tent of the testimony, and behold, the staff of Aaron for the house of Levi had sprouted and put forth buds and produced blossoms, and it bore ripe almonds.
NUM|17|9|Then Moses brought out all the staffs from before the LORD to all the people of Israel. And they looked, and each man took his staff.
NUM|17|10|And the LORD said to Moses, "Put back the staff of Aaron before the testimony, to be kept as a sign for the rebels, that you may make an end of their grumblings against me, lest they die."
NUM|17|11|Thus did Moses; as the LORD commanded him, so he did.
NUM|17|12|And the people of Israel said to Moses, "Behold, we perish, we are undone, we are all undone.
NUM|17|13|Everyone who comes near, who comes near to the tabernacle of the LORD, shall die. Are we all to perish?"
NUM|18|1|So the LORD said to Aaron, "You and your sons and your father's house with you shall bear iniquity connected with the sanctuary, and you and your sons with you shall bear iniquity connected with your priesthood.
NUM|18|2|And with you bring your brothers also, the tribe of Levi, the tribe of your father, that they may join you and minister to you while you and your sons with you are before the tent of the testimony.
NUM|18|3|They shall keep guard over you and over the whole tent, but shall not come near to the vessels of the sanctuary or to the altar lest they, and you, die.
NUM|18|4|They shall join you and keep guard over the tent of meeting for all the service of the tent, and no outsider shall come near you.
NUM|18|5|And you shall keep guard over the sanctuary and over the altar, that there may never again be wrath on the people of Israel.
NUM|18|6|And behold, I have taken your brothers the Levites from among the people of Israel. They are a gift to you, given to the LORD, to do the service of the tent of meeting.
NUM|18|7|And you and your sons with you shall guard your priesthood for all that concerns the altar and that is within the veil; and you shall serve. I give your priesthood as a gift, and any outsider who comes near shall be put to death."
NUM|18|8|Then the LORD spoke to Aaron, "Behold, I have given you charge of the contributions made to me, all the consecrated things of the people of Israel. I have given them to you as a portion and to your sons as a perpetual due.
NUM|18|9|This shall be yours of the most holy things, reserved from the fire: every offering of theirs, every grain offering of theirs and every sin offering of theirs and every guilt offering of theirs, which they render to me, shall be most holy to you and to your sons.
NUM|18|10|In a most holy place shall you eat it. Every male may eat it; it is holy to you.
NUM|18|11|This also is yours: the contribution of their gift, all the wave offerings of the people of Israel. I have given them to you, and to your sons and daughters with you, as a perpetual due. Everyone who is clean in your house may eat it.
NUM|18|12|All the best of the oil and all the best of the wine and of the grain, the firstfruits of what they give to the LORD, I give to you.
NUM|18|13|The first ripe fruits of all that is in their land, which they bring to the LORD, shall be yours. Everyone who is clean in your house may eat it.
NUM|18|14|Every devoted thing in Israel shall be yours.
NUM|18|15|Everything that opens the womb of all flesh, whether man or beast, which they offer to the LORD, shall be yours. Nevertheless, the firstborn of man you shall redeem, and the firstborn of unclean animals you shall redeem.
NUM|18|16|And their redemption price (at a month old you shall redeem them) you shall fix at five shekels in silver, according to the shekel of the sanctuary, which is twenty gerahs.
NUM|18|17|But the firstborn of a cow, or the firstborn of a sheep, or the firstborn of a goat, you shall not redeem; they are holy. You shall sprinkle their blood on the altar and shall burn their fat as a food offering, with a pleasing aroma to the LORD.
NUM|18|18|But their flesh shall be yours, as the breast that is waved and as the right thigh are yours.
NUM|18|19|All the holy contributions that the people of Israel present to the LORD I give to you, and to your sons and daughters with you, as a perpetual due. It is a covenant of salt forever before the LORD for you and for your offspring with you."
NUM|18|20|And the LORD said to Aaron, "You shall have no inheritance in their land, neither shall you have any portion among them. I am your portion and your inheritance among the people of Israel.
NUM|18|21|"To the Levites I have given every tithe in Israel for an inheritance, in return for their service that they do, their service in the tent of meeting,
NUM|18|22|so that the people of Israel do not come near the tent of meeting, lest they bear sin and die.
NUM|18|23|But the Levites shall do the service of the tent of meeting, and they shall bear their iniquity. It shall be a perpetual statute throughout your generations, and among the people of Israel they shall have no inheritance.
NUM|18|24|For the tithe of the people of Israel, which they present as a contribution to the LORD, I have given to the Levites for an inheritance. Therefore I have said of them that they shall have no inheritance among the people of Israel."
NUM|18|25|And the LORD spoke to Moses, saying,
NUM|18|26|"Moreover, you shall speak and say to the Levites, 'When you take from the people of Israel the tithe that I have given you from them for your inheritance, then you shall present a contribution from it to the LORD, a tithe of the tithe.
NUM|18|27|And your contribution shall be counted to you as though it were the grain of the threshing floor, and as the fullness of the winepress.
NUM|18|28|So you shall also present a contribution to the LORD from all your tithes, which you receive from the people of Israel. And from it you shall give the LORD's contribution to Aaron the priest.
NUM|18|29|Out of all the gifts to you, you shall present every contribution due to the LORD; from each its best part is to be dedicated.'
NUM|18|30|Therefore you shall say to them, 'When you have offered from it the best of it, then the rest shall be counted to the Levites as produce of the threshing floor, and as produce of the winepress.
NUM|18|31|And you may eat it in any place, you and your households, for it is your reward in return for your service in the tent of meeting.
NUM|18|32|And you shall bear no sin by reason of it, when you have contributed the best of it. But you shall not profane the holy things of the people of Israel, lest you die.'"
NUM|19|1|Now the LORD spoke to Moses and to Aaron, saying,
NUM|19|2|"This is the statute of the law that the LORD has commanded: Tell the people of Israel to bring you a red heifer without defect, in which there is no blemish, and on which a yoke has never come.
NUM|19|3|And you shall give it to Eleazar the priest, and it shall be taken outside the camp and slaughtered before him.
NUM|19|4|And Eleazar the priest shall take some of its blood with his finger, and sprinkle some of its blood toward the front of the tent of meeting seven times.
NUM|19|5|And the heifer shall be burned in his sight. Its skin, its flesh, and its blood, with its dung, shall be burned.
NUM|19|6|And the priest shall take cedarwood and hyssop and scarlet yarn, and throw them into the fire burning the heifer.
NUM|19|7|Then the priest shall wash his clothes and bathe his body in water, and afterward he may come into the camp. But the priest shall be unclean until evening.
NUM|19|8|The one who burns the heifer shall wash his clothes in water and bathe his body in water and shall be unclean until evening.
NUM|19|9|And a man who is clean shall gather up the ashes of the heifer and deposit them outside the camp in a clean place. And they shall be kept for the water for impurity for the congregation of the people of Israel; it is a sin offering.
NUM|19|10|And the one who gathers the ashes of the heifer shall wash his clothes and be unclean until evening. And this shall be a perpetual statute for the people of Israel, and for the stranger who sojourns among them.
NUM|19|11|"Whoever touches the dead body of any person shall be unclean seven days.
NUM|19|12|He shall cleanse himself with the water on the third day and on the seventh day, and so be clean. But if he does not cleanse himself on the third day and on the seventh day, he will not become clean.
NUM|19|13|Whoever touches a dead person, the body of anyone who has died, and does not cleanse himself, defiles the tabernacle of the LORD, and that person shall be cut off from Israel; because the water for impurity was not thrown on him, he shall be unclean. His uncleanness is still on him.
NUM|19|14|"This is the law when someone dies in a tent: everyone who comes into the tent and everyone who is in the tent shall be unclean seven days.
NUM|19|15|And every open vessel that has no cover fastened on it is unclean.
NUM|19|16|Whoever in the open field touches someone who was killed with a sword or who died naturally, or touches a human bone or a grave, shall be unclean seven days.
NUM|19|17|For the unclean they shall take some ashes of the burnt sin offering, and fresh water shall be added in a vessel.
NUM|19|18|Then a clean person shall take hyssop and dip it in the water and sprinkle it on the tent and on all the furnishings and on the persons who were there and on whoever touched the bone, or the slain or the dead or the grave.
NUM|19|19|And the clean person shall sprinkle it on the unclean on the third day and on the seventh day. Thus on the seventh day he shall cleanse him, and he shall wash his clothes and bathe himself in water, and at evening he shall be clean.
NUM|19|20|"If the man who is unclean does not cleanse himself, that person shall be cut off from the midst of the assembly, since he has defiled the sanctuary of the LORD. Because the water for impurity has not been thrown on him, he is unclean.
NUM|19|21|And it shall be a statute forever for them. The one who sprinkles the water for impurity shall wash his clothes, and the one who touches the water for impurity shall be unclean until evening.
NUM|19|22|And whatever the unclean person touches shall be unclean, and anyone who touches it shall be unclean until evening."
NUM|20|1|And the people of Israel, the whole congregation, came into the wilderness of Zin in the first month, and the people stayed in Kadesh. And Miriam died there and was buried there.
NUM|20|2|Now there was no water for the congregation. And they assembled themselves together against Moses and against Aaron.
NUM|20|3|And the people quarreled with Moses and said, "Would that we had perished when our brothers perished before the LORD!
NUM|20|4|Why have you brought the assembly of the LORD into this wilderness, that we should die here, both we and our cattle?
NUM|20|5|And why have you made us come up out of Egypt to bring us to this evil place? It is no place for grain or figs or vines or pomegranates, and there is no water to drink."
NUM|20|6|Then Moses and Aaron went from the presence of the assembly to the entrance of the tent of meeting and fell on their faces. And the glory of the LORD appeared to them,
NUM|20|7|and the LORD spoke to Moses, saying,
NUM|20|8|"Take the staff, and assemble the congregation, you and Aaron your brother, and tell the rock before their eyes to yield its water. So you shall bring water out of the rock for them and give drink to the congregation and their cattle."
NUM|20|9|And Moses took the staff from before the LORD, as he commanded him.
NUM|20|10|Then Moses and Aaron gathered the assembly together before the rock, and he said to them, "Hear now, you rebels: shall we bring water for you out of this rock?"
NUM|20|11|And Moses lifted up his hand and struck the rock with his staff twice, and water came out abundantly, and the congregation drank, and their livestock.
NUM|20|12|And the LORD said to Moses and Aaron, "Because you did not believe in me, to uphold me as holy in the eyes of the people of Israel, therefore you shall not bring this assembly into the land that I have given them."
NUM|20|13|These are the waters of Meribah, where the people of Israel quarreled with the LORD, and through them he showed himself holy.
NUM|20|14|Moses sent messengers from Kadesh to the king of Edom: "Thus says your brother Israel: You know all the hardship that we have met:
NUM|20|15|how our fathers went down to Egypt, and we lived in Egypt a long time. And the Egyptians dealt harshly with us and our fathers.
NUM|20|16|And when we cried to the LORD, he heard our voice and sent an angel and brought us out of Egypt. And here we are in Kadesh, a city on the edge of your territory.
NUM|20|17|Please let us pass through your land. We will not pass through field or vineyard, or drink water from a well. We will go along the King's Highway. We will not turn aside to the right hand or to the left until we have passed through your territory."
NUM|20|18|But Edom said to him, "You shall not pass through, lest I come out with the sword against you."
NUM|20|19|And the people of Israel said to him, "We will go up by the highway, and if we drink of your water, I and my livestock, then I will pay for it. Let me only pass through on foot, nothing more."
NUM|20|20|But he said, "You shall not pass through." And Edom came out against them with a large army and with a strong force.
NUM|20|21|Thus Edom refused to give Israel passage through his territory, so Israel turned away from him.
NUM|20|22|And they journeyed from Kadesh, and the people of Israel, the whole congregation, came to Mount Hor.
NUM|20|23|And the LORD said to Moses and Aaron at Mount Hor, on the border of the land of Edom,
NUM|20|24|"Let Aaron be gathered to his people, for he shall not enter the land that I have given to the people of Israel, because you rebelled against my command at the waters of Meribah.
NUM|20|25|Take Aaron and Eleazar his son and bring them up to Mount Hor.
NUM|20|26|And strip Aaron of his garments and put them on Eleazar his son. And Aaron shall be gathered to his people and shall die there."
NUM|20|27|Moses did as the LORD commanded. And they went up Mount Hor in the sight of all the congregation.
NUM|20|28|And Moses stripped Aaron of his garments and put them on Eleazar his son. And Aaron died there on the top of the mountain. Then Moses and Eleazar came down from the mountain.
NUM|20|29|And when all the congregation saw that Aaron had perished, all the house of Israel wept for Aaron thirty days.
NUM|21|1|When the Canaanite, the king of Arad, who lived in the Negeb, heard that Israel was coming by the way of Atharim, he fought against Israel, and took some of them captive.
NUM|21|2|And Israel vowed a vow to the LORD and said, "If you will indeed give this people into my hand, then I will devote their cities to destruction."
NUM|21|3|And the LORD obeyed the voice of Israel and gave over the Canaanites, and they devoted them and their cities to destruction. So the name of the place was called Hormah.
NUM|21|4|From Mount Hor they set out by the way to the Red Sea, to go around the land of Edom. And the people became impatient on the way.
NUM|21|5|And the people spoke against God and against Moses, "Why have you brought us up out of Egypt to die in the wilderness? For there is no food and no water, and we loathe this worthless food."
NUM|21|6|Then the LORD sent fiery serpents among the people, and they bit the people, so that many people of Israel died.
NUM|21|7|And the people came to Moses and said, "We have sinned, for we have spoken against the LORD and against you. Pray to the LORD, that he take away the serpents from us." So Moses prayed for the people.
NUM|21|8|And the LORD said to Moses, "Make a fiery serpent and set it on a pole, and everyone who is bitten, when he sees it, shall live."
NUM|21|9|So Moses made a bronze serpent and set it on a pole. And if a serpent bit anyone, he would look at the bronze serpent and live.
NUM|21|10|And the people of Israel set out and camped in Oboth.
NUM|21|11|And they set out from Oboth and camped at Iye-abarim, in the wilderness that is opposite Moab, toward the sunrise.
NUM|21|12|From there they set out and camped in the Valley of Zered.
NUM|21|13|From there they set out and camped on the other side of the Arnon, which is in the wilderness that extends from the border of the Amorites, for the Arnon is the border of Moab, between Moab and the Amorites.
NUM|21|14|Wherefore it is said in the Book of the Wars of the LORD, "Waheb in Suphah, and the valleys of the Arnon,
NUM|21|15|and the slope of the valleys that extends to the seat of Ar, and leans to the border of Moab."
NUM|21|16|And from there they continued to Beer; that is the well of which the LORD said to Moses, "Gather the people together, so that I may give them water."
NUM|21|17|Then Israel sang this song: "Spring up, O well!- Sing to it!-
NUM|21|18|the well that the princes dug, that the nobles of the people delved, with the scepter and with their staffs." And from the wilderness they went on to Mattanah,
NUM|21|19|and from Mattanah to Nahaliel, and from Nahaliel to Bamoth,
NUM|21|20|and from Bamoth to the valley lying in the region of Moab by the top of Pisgah that looks down on the desert.
NUM|21|21|Then Israel sent messengers to Sihon king of the Amorites, saying,
NUM|21|22|"Let me pass through your land. We will not turn aside into field or vineyard. We will not drink the water of a well. We will go by the King's Highway until we have passed through your territory."
NUM|21|23|But Sihon would not allow Israel to pass through his territory. He gathered all his people together and went out against Israel to the wilderness and came to Jahaz and fought against Israel.
NUM|21|24|And Israel defeated him with the edge of the sword and took possession of his land from the Arnon to the Jabbok, as far as to the Ammonites, for the border of the Ammonites was strong.
NUM|21|25|And Israel took all these cities, and Israel settled in all the cities of the Amorites, in Heshbon, and in all its villages.
NUM|21|26|For Heshbon was the city of Sihon the king of the Amorites, who had fought against the former king of Moab and taken all his land out of his hand, as far as the Arnon.
NUM|21|27|Therefore the ballad singers say, "Come to Heshbon, let it be built; let the city of Sihon be established.
NUM|21|28|For fire came out from Heshbon, flame from the city of Sihon. It devoured Ar of Moab, and swallowed the heights of the Arnon.
NUM|21|29|Woe to you, O Moab! You are undone, O people of Chemosh! He has made his sons fugitives, and his daughters captives, to an Amorite king, Sihon.
NUM|21|30|So we overthrew them; Heshbon, as far as Dibon, perished; and we laid waste as far as Nophah; fire spread as far as Medeba."
NUM|21|31|Thus Israel lived in the land of the Amorites.
NUM|21|32|And Moses sent to spy out Jazer, and they captured its villages and dispossessed the Amorites who were there.
NUM|21|33|Then they turned and went up by the way to Bashan. And Og the king of Bashan came out against them, he and all his people, to battle at Edrei.
NUM|21|34|But the LORD said to Moses, "Do not fear him, for I have given him into your hand, and all his people, and his land. And you shall do to him as you did to Sihon king of the Amorites, who lived at Heshbon."
NUM|21|35|So they defeated him and his sons and all his people, until he had no survivor left. And they possessed his land.
NUM|22|1|Then the people of Israel set out and camped in the plains of Moab beyond the Jordan at Jericho.
NUM|22|2|And Balak the son of Zippor saw all that Israel had done to the Amorites.
NUM|22|3|And Moab was in great dread of the people, because they were many. Moab was overcome with fear of the people of Israel.
NUM|22|4|And Moab said to the elders of Midian, "This horde will now lick up all that is around us, as the ox licks up the grass of the field." So Balak the son of Zippor, who was king of Moab at that time,
NUM|22|5|sent messengers to Balaam the son of Beor at Pethor, which is near the River in the land of the people of Amaw, to call him, saying, "Behold, a people has come out of Egypt. They cover the face of the earth, and they are dwelling opposite me.
NUM|22|6|Come now, curse this people for me, since they are too mighty for me. Perhaps I shall be able to defeat them and drive them from the land, for I know that he whom you bless is blessed, and he whom you curse is cursed."
NUM|22|7|So the elders of Moab and the elders of Midian departed with the fees for divination in their hand. And they came to Balaam and gave him Balak's message.
NUM|22|8|And he said to them, "Lodge here tonight, and I will bring back word to you, as the LORD speaks to me." So the princes of Moab stayed with Balaam.
NUM|22|9|And God came to Balaam and said, "Who are these men with you?"
NUM|22|10|And Balaam said to God, "Balak the son of Zippor, king of Moab, has sent to me, saying,
NUM|22|11|'Behold, a people has come out of Egypt, and it covers the face of the earth. Now come, curse them for me. Perhaps I shall be able to fight against them and drive them out.'"
NUM|22|12|God said to Balaam, "You shall not go with them. You shall not curse the people, for they are blessed."
NUM|22|13|So Balaam rose in the morning and said to the princes of Balak, "Go to your own land, for the LORD has refused to let me go with you."
NUM|22|14|So the princes of Moab rose and went to Balak and said, "Balaam refuses to come with us."
NUM|22|15|Once again Balak sent princes, more in number and more honorable than these.
NUM|22|16|And they came to Balaam and said to him, "Thus says Balak the son of Zippor: 'Let nothing hinder you from coming to me,
NUM|22|17|for I will surely do you great honor, and whatever you say to me I will do. Come, curse this people for me.'"
NUM|22|18|But Balaam answered and said to the servants of Balak, "Though Balak were to give me his house full of silver and gold, I could not go beyond the command of the LORD my God to do less or more.
NUM|22|19|So you, too, please stay here tonight, that I may know what more the LORD will say to me."
NUM|22|20|And God came to Balaam at night and said to him, "If the men have come to call you, rise, go with them; but only do what I tell you."
NUM|22|21|So Balaam rose in the morning and saddled his donkey and went with the princes of Moab.
NUM|22|22|But God's anger was kindled because he went, and the angel of the LORD took his stand in the way as his adversary. Now he was riding on the donkey, and his two servants were with him.
NUM|22|23|And the donkey saw the angel of the LORD standing in the road, with a drawn sword in his hand. And the donkey turned aside out of the road and went into the field. And Balaam struck the donkey, to turn her into the road.
NUM|22|24|Then the angel of the LORD stood in a narrow path between the vineyards, with a wall on either side.
NUM|22|25|And when the donkey saw the angel of the LORD, she pushed against the wall and pressed Balaam's foot against the wall. So he struck her again.
NUM|22|26|Then the angel of the LORD went ahead and stood in a narrow place, where there was no way to turn either to the right or to the left.
NUM|22|27|When the donkey saw the angel of the LORD, she lay down under Balaam. And Balaam's anger was kindled, and he struck the donkey with his staff.
NUM|22|28|Then the LORD opened the mouth of the donkey, and she said to Balaam, "What have I done to you, that you have struck me these three times?"
NUM|22|29|And Balaam said to the donkey, "Because you have made a fool of me. I wish I had a sword in my hand, for then I would kill you."
NUM|22|30|And the donkey said to Balaam, "Am I not your donkey, on which you have ridden all your life long to this day? Is it my habit to treat you this way?" And he said, "No."
NUM|22|31|Then the LORD opened the eyes of Balaam, and he saw the angel of the LORD standing in the way, with his drawn sword in his hand. And he bowed down and fell on his face.
NUM|22|32|And the angel of the LORD said to him, "Why have you struck your donkey these three times? Behold, I have come out to oppose you because your way is perverse before me.
NUM|22|33|The donkey saw me and turned aside before me these three times. If she had not turned aside from me, surely just now I would have killed you and let her live."
NUM|22|34|Then Balaam said to the angel of the LORD, "I have sinned, for I did not know that you stood in the road against me. Now therefore, if it is evil in your sight, I will turn back."
NUM|22|35|And the angel of the LORD said to Balaam, "Go with the men, but speak only the word that I tell you." So Balaam went on with the princes of Balak.
NUM|22|36|When Balak heard that Balaam had come, he went out to meet him at the city of Moab, on the border formed by the Arnon, at the extremity of the border.
NUM|22|37|And Balak said to Balaam, "Did I not send to you to call you? Why did you not come to me? Am I not able to honor you?"
NUM|22|38|Balaam said to Balak, "Behold, I have come to you! Have I now any power of my own to speak anything? The word that God puts in my mouth, that must I speak."
NUM|22|39|Then Balaam went with Balak, and they came to Kiriath-huzoth.
NUM|22|40|And Balak sacrificed oxen and sheep, and sent for Balaam and for the princes who were with him.
NUM|22|41|And in the morning Balak took Balaam and brought him up to Bamoth-baal, and from there he saw a fraction of the people.
NUM|23|1|And Balaam said to Balak, "Build for me here seven altars, and prepare for me here seven bulls and seven rams."
NUM|23|2|Balak did as Balaam had said. And Balak and Balaam offered on each altar a bull and a ram.
NUM|23|3|And Balaam said to Balak, "Stand beside your burnt offering, and I will go. Perhaps the LORD will come to meet me, and whatever he shows me I will tell you." And he went to a bare height,
NUM|23|4|and God met Balaam. And Balaam said to him, "I have arranged the seven altars and I have offered on each altar a bull and a ram."
NUM|23|5|And the LORD put a word in Balaam's mouth and said, "Return to Balak, and thus you shall speak."
NUM|23|6|And he returned to him, and behold, he and all the princes of Moab were standing beside his burnt offering.
NUM|23|7|And Balaam took up his discourse and said, "From Aram Balak has brought me, the king of Moab from the eastern mountains: 'Come, curse Jacob for me, and come, denounce Israel!'
NUM|23|8|How can I curse whom God has not cursed? How can I denounce whom the LORD has not denounced?
NUM|23|9|For from the top of the crags I see him, from the hills I behold him; behold, a people dwelling alone, and not counting itself among the nations!
NUM|23|10|Who can count the dust of Jacob or number the fourth part of Israel? Let me die the death of the upright, and let my end be like his!"
NUM|23|11|And Balak said to Balaam, "What have you done to me? I took you to curse my enemies, and behold, you have done nothing but bless them."
NUM|23|12|And he answered and said, "Must I not take care to speak what the LORD puts in my mouth?"
NUM|23|13|And Balak said to him, "Please come with me to another place, from which you may see them. You shall see only a fraction of them and shall not see them all. Then curse them for me from there."
NUM|23|14|And he took him to the field of Zophim, to the top of Pisgah, and built seven altars and offered a bull and a ram on each altar.
NUM|23|15|Balaam said to Balak, "Stand here beside your burnt offering, while I meet the LORD over there."
NUM|23|16|And the LORD met Balaam and put a word in his mouth and said, "Return to Balak, and thus shall you speak."
NUM|23|17|And he came to him, and behold, he was standing beside his burnt offering, and the princes of Moab with him. And Balak said to him, "What has the LORD spoken?"
NUM|23|18|And Balaam took up his discourse and said, "Rise, Balak, and hear; give ear to me, O son of Zippor:
NUM|23|19|God is not man, that he should lie, or a son of man, that he should change his mind. Has he said, and will he not do it? Or has he spoken, and will he not fulfill it?
NUM|23|20|Behold, I received a command to bless: he has blessed, and I cannot revoke it.
NUM|23|21|He has not beheld misfortune in Jacob, nor has he seen trouble in Israel. The LORD their God is with them, and the shout of a king is among them.
NUM|23|22|God brings them out of Egypt and is for them like the horns of the wild ox.
NUM|23|23|For there is no enchantment against Jacob, no divination against Israel; now it shall be said of Jacob and Israel, 'What has God wrought!'
NUM|23|24|Behold, a people! As a lioness it rises up and as a lion it lifts itself; it does not lie down until it has devoured the prey and drunk the blood of the slain."
NUM|23|25|And Balak said to Balaam, "Do not curse them at all, and do not bless them at all."
NUM|23|26|But Balaam answered Balak, "Did I not tell you, 'All that the LORD says, that I must do'?"
NUM|23|27|And Balak said to Balaam, "Come now, I will take you to another place. Perhaps it will please God that you may curse them for me from there."
NUM|23|28|So Balak took Balaam to the top of Peor, which overlooks the desert.
NUM|23|29|And Balaam said to Balak, "Build for me here seven altars and prepare for me here seven bulls and seven rams."
NUM|23|30|And Balak did as Balaam had said, and offered a bull and a ram on each altar.
NUM|24|1|When Balaam saw that it pleased the LORD to bless Israel, he did not go, as at other times, to look for omens, but set his face toward the wilderness.
NUM|24|2|And Balaam lifted up his eyes and saw Israel camping tribe by tribe. And the Spirit of God came upon him,
NUM|24|3|and he took up his discourse and said, "The oracle of Balaam the son of Beor, the oracle of the man whose eye is opened,
NUM|24|4|the oracle of him who hears the words of God, who sees the vision of the Almighty, falling down with his eyes uncovered:
NUM|24|5|How lovely are your tents, O Jacob, your encampments, O Israel!
NUM|24|6|Like palm groves that stretch afar, like gardens beside a river, like aloes that the LORD has planted, like cedar trees beside the waters.
NUM|24|7|Water shall flow from his buckets, and his seed shall be in many waters; his king shall be higher than Agag, and his kingdom shall be exalted.
NUM|24|8|God brings him out of Egypt and is for him like the horns of the wild ox; he shall eat up the nations, his adversaries, and shall break their bones in pieces and pierce them through with his arrows.
NUM|24|9|He crouched, he lay down like a lion and like a lioness; who will rouse him up? Blessed are those who bless you, and cursed are those who curse you."
NUM|24|10|And Balak's anger was kindled against Balaam, and he struck his hands together. And Balak said to Balaam, "I called you to curse my enemies, and behold, you have blessed them these three times.
NUM|24|11|Therefore now flee to your own place. I said, 'I will certainly honor you,' but the LORD has held you back from honor."
NUM|24|12|And Balaam said to Balak, "Did I not tell your messengers whom you sent to me,
NUM|24|13|'If Balak should give me his house full of silver and gold, I would not be able to go beyond the word of the LORD, to do either good or bad of my own will. What the LORD speaks, that will I speak'?
NUM|24|14|And now, behold, I am going to my people. Come, I will let you know what this people will do to your people in the latter days."
NUM|24|15|And he took up his discourse and said, "The oracle of Balaam the son of Beor, the oracle of the man whose eye is opened,
NUM|24|16|the oracle of him who hears the words of God, and knows the knowledge of the Most High, who sees the vision of the Almighty, falling down with his eyes uncovered:
NUM|24|17|I see him, but not now; I behold him, but not near: a star shall come out of Jacob, and a scepter shall rise out of Israel; it shall crush the forehead of Moab and break down all the sons of Sheth.
NUM|24|18|Edom shall be dispossessed; Seir also, his enemies, shall be dispossessed. Israel is doing valiantly.
NUM|24|19|And one from Jacob shall exercise dominion and destroy the survivors of cities!"
NUM|24|20|Then he looked on Amalek and took up his discourse and said, "Amalek was the first among the nations, but its end is utter destruction."
NUM|24|21|And he looked on the Kenite, and took up his discourse and said, "Enduring is your dwelling place, and your nest is set in the rock.
NUM|24|22|Nevertheless, Kain shall be burned when Asshur takes you away captive."
NUM|24|23|And he took up his discourse and said, "Alas, who shall live when God does this?
NUM|24|24|But ships shall come from Kittim and shall afflict Asshur and Eber; and he too shall come to utter destruction."
NUM|24|25|Then Balaam rose and went back to his place. And Balak also went his way.
NUM|25|1|While Israel lived in Shittim, the people began to whore with the daughters of Moab.
NUM|25|2|These invited the people to the sacrifices of their gods, and the people ate and bowed down to their gods.
NUM|25|3|So Israel yoked himself to Baal of Peor. And the anger of the LORD was kindled against Israel.
NUM|25|4|And the LORD said to Moses, "Take all the chiefs of the people and hang them in the sun before the LORD, that the fierce anger of the LORD may turn away from Israel."
NUM|25|5|And Moses said to the judges of Israel, "Each of you kill those of his men who have yoked themselves to Baal of Peor."
NUM|25|6|And behold, one of the people of Israel came and brought a Midianite woman to his family, in the sight of Moses and in the sight of the whole congregation of the people of Israel, while they were weeping in the entrance of the tent of meeting.
NUM|25|7|When Phinehas the son of Eleazar, son of Aaron the priest, saw it, he rose and left the congregation and took a spear in his hand
NUM|25|8|and went after the man of Israel into the chamber and pierced both of them, the man of Israel and the woman through her belly. Thus the plague on the people of Israel was stopped.
NUM|25|9|Nevertheless, those who died by the plague were twenty-four thousand.
NUM|25|10|And the LORD said to Moses,
NUM|25|11|"Phinehas the son of Eleazar, son of Aaron the priest, has turned back my wrath from the people of Israel, in that he was jealous with my jealousy among them, so that I did not consume the people of Israel in my jealousy.
NUM|25|12|Therefore say, 'Behold, I give to him my covenant of peace,
NUM|25|13|and it shall be to him and to his descendants after him the covenant of a perpetual priesthood, because he was jealous for his God and made atonement for the people of Israel.'"
NUM|25|14|The name of the slain man of Israel, who was killed with the Midianite woman, was Zimri the son of Salu, chief of a father's house belonging to the Simeonites.
NUM|25|15|And the name of the Midianite woman who was killed was Cozbi the daughter of Zur, who was the tribal head of a father's house in Midian.
NUM|25|16|And the LORD spoke to Moses, saying,
NUM|25|17|"Harass the Midianites and strike them down,
NUM|25|18|for they have harassed you with their wiles, with which they beguiled you in the matter of Peor, and in the matter of Cozbi, the daughter of the chief of Midian, their sister, who was killed on the day of the plague on account of Peor."
NUM|26|1|After the plague, the LORD said to Moses and to Eleazar the son of Aaron, the priest,
NUM|26|2|"Take a census of all the congregation of the people of Israel, from twenty years old and upward, by their fathers' houses, all in Israel who are able to go to war."
NUM|26|3|And Moses and Eleazar the priest spoke with them in the plains of Moab by the Jordan at Jericho, saying,
NUM|26|4|"Take a census of the people, from twenty years old and upward," as the LORD commanded Moses. The people of Israel who came out of the land of Egypt were:
NUM|26|5|Reuben, the firstborn of Israel; the sons of Reuben: of Hanoch, the clan of the Hanochites; of Pallu, the clan of the Palluites;
NUM|26|6|of Hezron, the clan of the Hezronites; of Carmi, the clan of the Carmites.
NUM|26|7|These are the clans of the Reubenites, and those listed were 43,730.
NUM|26|8|And the sons of Pallu: Eliab.
NUM|26|9|The sons of Eliab: Nemuel, Dathan, and Abiram. These are the Dathan and Abiram, chosen from the congregation, who contended against Moses and Aaron in the company of Korah, when they contended against the LORD
NUM|26|10|and the earth opened its mouth and swallowed them up together with Korah, when that company died, when the fire devoured 250 men, and they became a warning.
NUM|26|11|But the sons of Korah did not die.
NUM|26|12|The sons of Simeon according to their clans: of Nemuel, the clan of the Nemuelites; of Jamin, the clan of the Ja-minites; of Jachin, the clan of the Jachinites;
NUM|26|13|of Zerah, the clan of the Zerahites; of Shaul, the clan of the Sha-ulites.
NUM|26|14|These are the clans of the Simeonites, 22,200.
NUM|26|15|The sons of Gad according to their clans: of Zephon, the clan of the Zephonites; of Haggi, the clan of the Haggites; of Shuni, the clan of the Shunites;
NUM|26|16|of Ozni, the clan of the Oznites; of Eri, the clan of the Erites;
NUM|26|17|of Arod, the clan of the Arodites; of Areli, the clan of the Arelites.
NUM|26|18|These are the clans of the sons of Gad as they were listed, 40,500.
NUM|26|19|The sons of Judah were Er and Onan; and Er and Onan died in the land of Canaan.
NUM|26|20|And the sons of Judah according to their clans were: of Shelah, the clan of the Shelanites; of Perez, the clan of the Perezites; of Zerah, the clan of the Zerahites.
NUM|26|21|And the sons of Perez were: of Hezron, the clan of the Hezronites; of Hamul, the clan of the Hamulites.
NUM|26|22|These are the clans of Judah as they were listed, 76,500.
NUM|26|23|The sons of Issachar according to their clans: of Tola, the clan of the Tolaites; of Puvah, the clan of the Punites;
NUM|26|24|of Jashub, the clan of the Ja-shubites; of Shimron, the clan of the Shimronites.
NUM|26|25|These are the clans of Issachar as they were listed, 64,300.
NUM|26|26|The sons of Zebulun, according to their clans: of Sered, the clan of the Seredites; of Elon, the clan of the Elonites; of Jahleel, the clan of the Jah-leelites.
NUM|26|27|These are the clans of the Zeb-ulunites as they were listed, 60,500.
NUM|26|28|The sons of Joseph according to their clans: Manasseh and Ephraim.
NUM|26|29|The sons of Manasseh: of Machir, the clan of the Machirites; and Machir was the father of Gilead; of Gilead, the clan of the Gileadites.
NUM|26|30|These are the sons of Gilead: of Iezer, the clan of the Iezerites; of Helek, the clan of the Helekites;
NUM|26|31|and of Asriel, the clan of the Asrielites; and of Shechem, the clan of the Shechemites;
NUM|26|32|and of Shemida, the clan of the Shemidaites; and of Hepher, the clan of the Hepherites.
NUM|26|33|Now Zelophehad the son of Hepher had no sons, but daughters. And the names of the daughters of Zelophehad were Mahlah, Noah, Hoglah, Milcah, and Tirzah.
NUM|26|34|These are the clans of Manasseh, and those listed were 52,700.
NUM|26|35|These are the sons of Ephraim according to their clans: of Shuthelah, the clan of the Shuthelahites; of Becher, the clan of the Becherites; of Tahan, the clan of the Tahanites.
NUM|26|36|And these are the sons of Shuthelah: of Eran, the clan of the Eranites.
NUM|26|37|These are the clans of the sons of Ephraim as they were listed, 32,500. These are the sons of Joseph according to their clans.
NUM|26|38|The sons of Benjamin according to their clans: of Bela, the clan of the Belaites; of Ashbel, the clan of the Ashbelites; of Ahiram, the clan of the Ahiramites;
NUM|26|39|of Shephupham, the clan of the Shuphamites; of Hupham, the clan of the Huphamites.
NUM|26|40|And the sons of Bela were Ard and Naaman: of Ard, the clan of the Ardites; of Naaman, the clan of the Naamites.
NUM|26|41|These are the sons of Benjamin according to their clans, and those listed were 45,600.
NUM|26|42|These are the sons of Dan according to their clans: of Shuham, the clan of the Shuhamites. These are the clans of Dan according to their clans.
NUM|26|43|All the clans of the Shuhamites, as they were listed, were 64,400.
NUM|26|44|The sons of Asher according to their clans: of Imnah, the clan of the Imnites; of Ishvi, the clan of the Ishvites; of Beriah, the clan of the Beriites.
NUM|26|45|Of the sons of Beriah: of Heber, the clan of the Heberites; of Malchiel, the clan of the Malchielites.
NUM|26|46|And the name of the daughter of Asher was Serah.
NUM|26|47|These are the clans of the sons of Asher as they were listed, 53,400.
NUM|26|48|The sons of Naphtali according to their clans: of Jahzeel, the clan of the Jahzeelites; of Guni, the clan of the Gunites;
NUM|26|49|of Jezer, the clan of the Jezerites; of Shillem, the clan of the Shillemites.
NUM|26|50|These are the clans of Naphtali according to their clans, and those listed were 45,400.
NUM|26|51|This was the list of the people of Israel, 601,730.
NUM|26|52|The LORD spoke to Moses, saying,
NUM|26|53|"Among these the land shall be divided for inheritance according to the number of names.
NUM|26|54|To a large tribe you shall give a large inheritance, and to a small tribe you shall give a small inheritance; every tribe shall be given its inheritance in proportion to its list.
NUM|26|55|But the land shall be divided by lot. According to the names of the tribes of their fathers they shall inherit.
NUM|26|56|Their inheritance shall be divided according to lot between the larger and the smaller."
NUM|26|57|This was the list of the Levites according to their clans: of Gershon, the clan of the Gershonites; of Kohath, the clan of the Kohathites; of Merari, the clan of the Merarites.
NUM|26|58|These are the clans of Levi: the clan of the Libnites, the clan of the Hebronites, the clan of the Mahlites, the clan of the Mushites, the clan of the Korahites. And Kohath was the father of Amram.
NUM|26|59|The name of Amram's wife was Jochebed the daughter of Levi, who was born to Levi in Egypt. And she bore to Amram Aaron and Moses and Miriam their sister.
NUM|26|60|And to Aaron were born Nadab, Abihu, Eleazar, and Ithamar.
NUM|26|61|But Nadab and Abihu died when they offered unauthorized fire before the LORD.
NUM|26|62|And those listed were 23,000, every male from a month old and upward. For they were not listed among the people of Israel, because there was no inheritance given to them among the people of Israel.
NUM|26|63|These were those listed by Moses and Eleazar the priest, who listed the people of Israel in the plains of Moab by the Jordan at Jericho.
NUM|26|64|But among these there was not one of those listed by Moses and Aaron the priest, who had listed the people of Israel in the wilderness of Sinai.
NUM|26|65|For the LORD had said of them, "They shall die in the wilderness." Not one of them was left, except Caleb the son of Jephunneh and Joshua the son of Nun.
NUM|27|1|Then drew near the daughters of Zelophehad the son of Hepher, son of Gilead, son of Machir, son of Manasseh, from the clans of Manasseh the son of Joseph. The names of his daughters were: Mahlah, Noah, Hoglah, Milcah, and Tirzah.
NUM|27|2|And they stood before Moses and before Eleazar the priest and before the chiefs and all the congregation, at the entrance of the tent of meeting, saying,
NUM|27|3|"Our father died in the wilderness. He was not among the company of those who gathered themselves together against the LORD in the company of Korah, but died for his own sin. And he had no sons.
NUM|27|4|Why should the name of our father be taken away from his clan because he had no son? Give to us a possession among our father's brothers."
NUM|27|5|Moses brought their case before the LORD.
NUM|27|6|And the LORD said to Moses,
NUM|27|7|"The daughters of Zelophehad are right. You shall give them possession of an inheritance among their father's brothers and transfer the inheritance of their father to them.
NUM|27|8|And you shall speak to the people of Israel, saying, 'If a man dies and has no son, then you shall transfer his inheritance to his daughter.
NUM|27|9|And if he has no daughter, then you shall give his inheritance to his brothers.
NUM|27|10|And if he has no brothers, then you shall give his inheritance to his father's brothers.
NUM|27|11|And if his father has no brothers, then you shall give his inheritance to the nearest kinsman of his clan, and he shall possess it. And it shall be for the people of Israel a statute and rule, as the LORD commanded Moses.'"
NUM|27|12|The LORD said to Moses, "Go up into this mountain of Abarim and see the land that I have given to the people of Israel.
NUM|27|13|When you have seen it, you also shall be gathered to your people, as your brother Aaron was,
NUM|27|14|because you rebelled against my word in the wilderness of Zin when the congregation quarreled, failing to uphold me as holy at the waters before their eyes." (These are the waters of Meribah of Kadesh in the wilderness of Zin.)
NUM|27|15|Moses spoke to the LORD, saying,
NUM|27|16|"Let the LORD, the God of the spirits of all flesh, appoint a man over the congregation
NUM|27|17|who shall go out before them and come in before them, who shall lead them out and bring them in, that the congregation of the LORD may not be as sheep that have no shepherd."
NUM|27|18|So the LORD said to Moses, "Take Joshua the son of Nun, a man in whom is the Spirit, and lay your hand on him.
NUM|27|19|Make him stand before Eleazar the priest and all the congregation, and you shall commission him in their sight.
NUM|27|20|You shall invest him with some of your authority, that all the congregation of the people of Israel may obey.
NUM|27|21|And he shall stand before Eleazar the priest, who shall inquire for him by the judgment of the Urim before the LORD. At his word they shall go out, and at his word they shall come in, both he and all the people of Israel with him, the whole congregation."
NUM|27|22|And Moses did as the LORD commanded him. He took Joshua and made him stand before Eleazar the priest and the whole congregation,
NUM|27|23|and he laid his hands on him and commissioned him as the LORD directed through Moses.
NUM|28|1|The LORD spoke to Moses, saying,
NUM|28|2|"Command the people of Israel and say to them, 'My offering, my food for my food offerings, my pleasing aroma, you shall be careful to offer to me at its appointed time.'
NUM|28|3|And you shall say to them, This is the food offering that you shall offer to the LORD: two male lambs a year old without blemish, day by day, as a regular offering.
NUM|28|4|The one lamb you shall offer in the morning, and the other lamb you shall offer at twilight;
NUM|28|5|also a tenth of an ephah of fine flour for a grain offering, mixed with a quarter of a hin of beaten oil.
NUM|28|6|It is a regular burnt offering, which was ordained at Mount Sinai for a pleasing aroma, a food offering to the LORD.
NUM|28|7|Its drink offering shall be a quarter of a hin for each lamb. In the Holy Place you shall pour out a drink offering of strong drink to the LORD.
NUM|28|8|The other lamb you shall offer at twilight. Like the grain offering of the morning, and like its drink offering, you shall offer it as a food offering, with a pleasing aroma to the LORD.
NUM|28|9|"On the Sabbath day, two male lambs a year old without blemish, and two tenths of an ephah of fine flour for a grain offering, mixed with oil, and its drink offering:
NUM|28|10|this is the burnt offering of every Sabbath, besides the regular burnt offering and its drink offering.
NUM|28|11|"At the beginnings of your months, you shall offer a burnt offering to the LORD: two bulls from the herd, one ram, seven male lambs a year old without blemish;
NUM|28|12|also three tenths of an ephah of fine flour for a grain offering, mixed with oil, for each bull, and two tenths of fine flour for a grain offering, mixed with oil, for the one ram;
NUM|28|13|and a tenth of fine flour mixed with oil as a grain offering for every lamb; for a burnt offering with a pleasing aroma, a food offering to the LORD.
NUM|28|14|Their drink offerings shall be half a hin of wine for a bull, a third of a hin for a ram, and a quarter of a hin for a lamb. This is the burnt offering of each month throughout the months of the year.
NUM|28|15|Also one male goat for a sin offering to the LORD; it shall be offered besides the regular burnt offering and its drink offering.
NUM|28|16|"On the fourteenth day of the first month is the LORD's Passover,
NUM|28|17|and on the fifteenth day of this month is a feast. Seven days shall unleavened bread be eaten.
NUM|28|18|On the first day there shall be a holy convocation. You shall not do any ordinary work,
NUM|28|19|but offer a food offering, a burnt offering to the LORD: two bulls from the herd, one ram, and seven male lambs a year old; see that they are without blemish;
NUM|28|20|also their grain offering of fine flour mixed with oil; three tenths of an ephah shall you offer for a bull, and two tenths for a ram;
NUM|28|21|a tenth shall you offer for each of the seven lambs;
NUM|28|22|also one male goat for a sin offering, to make atonement for you.
NUM|28|23|You shall offer these besides the burnt offering of the morning, which is for a regular burnt offering.
NUM|28|24|In the same way you shall offer daily, for seven days, the food of a food offering, with a pleasing aroma to the LORD. It shall be offered besides the regular burnt offering and its drink offering.
NUM|28|25|And on the seventh day you shall have a holy convocation. You shall not do any ordinary work.
NUM|28|26|"On the day of the firstfruits, when you offer a grain offering of new grain to the LORD at your Feast of Weeks, you shall have a holy convocation. You shall not do any ordinary work,
NUM|28|27|but offer a burnt offering, with a pleasing aroma to the LORD: two bulls from the herd, one ram, seven male lambs a year old;
NUM|28|28|also their grain offering of fine flour mixed with oil, three tenths of an ephah for each bull, two tenths for one ram,
NUM|28|29|a tenth for each of the seven lambs;
NUM|28|30|with one male goat, to make atonement for you.
NUM|28|31|Besides the regular burnt offering and its grain offering, you shall offer them and their drink offering. See that they are without blemish.
NUM|29|1|"On the first day of the seventh month you shall have a holy convocation. You shall not do any ordinary work. It is a day for you to blow the trumpets,
NUM|29|2|and you shall offer a burnt offering, for a pleasing aroma to the LORD: one bull from the herd, one ram, seven male lambs a year old without blemish;
NUM|29|3|also their grain offering of fine flour mixed with oil, three tenths of an ephah for the bull, two tenths for the ram,
NUM|29|4|and one tenth for each of the seven lambs;
NUM|29|5|with one male goat for a sin offering, to make atonement for you;
NUM|29|6|besides the burnt offering of the new moon, and its grain offering, and the regular burnt offering and its grain offering, and their drink offering, according to the rule for them, for a pleasing aroma, a food offering to the LORD.
NUM|29|7|"On the tenth day of this seventh month you shall have a holy convocation and afflict yourselves. You shall do no work,
NUM|29|8|but you shall offer a burnt offering to the LORD, a pleasing aroma: one bull from the herd, one ram, seven male lambs a year old: see that they are without blemish.
NUM|29|9|And their grain offering shall be of fine flour mixed with oil, three tenths of an ephah for the bull, two tenths for the one ram,
NUM|29|10|a tenth for each of the seven lambs:
NUM|29|11|also one male goat for a sin offering, besides the sin offering of atonement, and the regular burnt offering and its grain offering, and their drink offerings.
NUM|29|12|"On the fifteenth day of the seventh month you shall have a holy convocation. You shall not do any ordinary work, and you shall keep a feast to the LORD seven days.
NUM|29|13|And you shall offer a burnt offering, a food offering, with a pleasing aroma to the LORD, thirteen bulls from the herd, two rams, fourteen male lambs a year old; they shall be without blemish;
NUM|29|14|and their grain offering of fine flour mixed with oil, three tenths of an ephah for each of the thirteen bulls, two tenths for each of the two rams,
NUM|29|15|and a tenth for each of the fourteen lambs;
NUM|29|16|also one male goat for a sin offering, besides the regular burnt offering, its grain offering and its drink offering.
NUM|29|17|"On the second day twelve bulls from the herd, two rams, fourteen male lambs a year old without blemish,
NUM|29|18|with the grain offering and the drink offerings for the bulls, for the rams, and for the lambs, in the prescribed quantities;
NUM|29|19|also one male goat for a sin offering, besides the regular burnt offering and its grain offering, and their drink offerings.
NUM|29|20|"On the third day eleven bulls, two rams, fourteen male lambs a year old without blemish,
NUM|29|21|with the grain offering and the drink offerings for the bulls, for the rams, and for the lambs, in the prescribed quantities;
NUM|29|22|also one male goat for a sin offering, besides the regular burnt offering and its grain offering and its drink offering.
NUM|29|23|"On the fourth day ten bulls, two rams, fourteen male lambs a year old without blemish,
NUM|29|24|with the grain offering and the drink offerings for the bulls, for the rams, and for the lambs, in the prescribed quantities;
NUM|29|25|also one male goat for a sin offering, besides the regular burnt offering, its grain offering and its drink offering.
NUM|29|26|"On the fifth day nine bulls, two rams, fourteen male lambs a year old without blemish,
NUM|29|27|with the grain offering and the drink offerings for the bulls, for the rams, and for the lambs, in the prescribed quantities;
NUM|29|28|also one male goat for a sin offering; besides the regular burnt offering and its grain offering and its drink offering.
NUM|29|29|"On the sixth day eight bulls, two rams, fourteen male lambs a year old without blemish,
NUM|29|30|with the grain offering and the drink offerings for the bulls, for the rams, and for the lambs, in the prescribed quantities;
NUM|29|31|also one male goat for a sin offering; besides the regular burnt offering, its grain offering, and its drink offerings.
NUM|29|32|"On the seventh day seven bulls, two rams, fourteen male lambs a year old without blemish,
NUM|29|33|with the grain offering and the drink offerings for the bulls, for the rams, and for the lambs, in the prescribed quantities;
NUM|29|34|also one male goat for a sin offering; besides the regular burnt offering, its grain offering, and its drink offering.
NUM|29|35|"On the eighth day you shall have a solemn assembly. You shall not do any ordinary work,
NUM|29|36|but you shall offer a burnt offering, a food offering, with a pleasing aroma to the LORD: one bull, one ram, seven male lambs a year old without blemish,
NUM|29|37|and the grain offering and the drink offerings for the bull, for the ram, and for the lambs, in the prescribed quantities;
NUM|29|38|also one male goat for a sin offering; besides the regular burnt offering and its grain offering and its drink offering.
NUM|29|39|"These you shall offer to the LORD at your appointed feasts, in addition to your vow offerings and your freewill offerings, for your burnt offerings, and for your grain offerings, and for your drink offerings, and for your peace offerings."
NUM|29|40|So Moses told the people of Israel everything just as the LORD had commanded Moses.
NUM|30|1|Moses spoke to the heads of the tribes of the people of Israel, saying, "This is what the LORD has commanded.
NUM|30|2|If a man vows a vow to the LORD, or swears an oath to bind himself by a pledge, he shall not break his word. He shall do according to all that proceeds out of his mouth.
NUM|30|3|If a woman vows a vow to the LORD and binds herself by a pledge, while within her father's house in her youth,
NUM|30|4|and her father hears of her vow and of her pledge by which she has bound herself and says nothing to her, then all her vows shall stand, and every pledge by which she has bound herself shall stand.
NUM|30|5|But if her father opposes her on the day that he hears of it, no vow of hers, no pledge by which she has bound herself shall stand. And the LORD will forgive her, because her father opposed her.
NUM|30|6|If she marries a husband, while under her vows or any thoughtless utterance of her lips by which she has bound herself,
NUM|30|7|and her husband hears of it and says nothing to her on the day that he hears, then her vows shall stand, and her pledges by which she has bound herself shall stand.
NUM|30|8|But if, on the day that her husband comes to hear of it, he opposes her, then he makes void her vow that was on her, and the thoughtless utterance of her lips by which she bound herself. And the LORD will forgive her.
NUM|30|9|(But any vow of a widow or of a divorced woman, anything by which she has bound herself, shall stand against her.)
NUM|30|10|And if she vowed in her husband's house or bound herself by a pledge with an oath,
NUM|30|11|and her husband heard of it and said nothing to her and did not oppose her, then all her vows shall stand, and every pledge by which she bound herself shall stand.
NUM|30|12|But if her husband makes them null and void on the day that he hears them, then whatever proceeds out of her lips concerning her vows or concerning her pledge of herself shall not stand. Her husband has made them void, and the LORD will forgive her.
NUM|30|13|Any vow and any binding oath to afflict herself, her husband may establish, or her husband may make void.
NUM|30|14|But if her husband says nothing to her from day to day, then he establishes all her vows or all her pledges that are upon her. He has established them, because he said nothing to her on the day that he heard of them.
NUM|30|15|But if he makes them null and void after he has heard of them, then he shall bear her iniquity."
NUM|30|16|These are the statutes that the LORD commanded Moses about a man and his wife and about a father and his daughter while she is in her youth within her father's house.
NUM|31|1|The LORD spoke to Moses, saying,
NUM|31|2|"Avenge the people of Israel on the Midianites. Afterward you shall be gathered to your people."
NUM|31|3|So Moses spoke to the people, saying, "Arm men from among you for the war, that they may go against Midian to execute the LORD's vengeance on Midian.
NUM|31|4|You shall send a thousand from each of the tribes of Israel to the war."
NUM|31|5|So there were provided, out of the thousands of Israel, a thousand from each tribe, twelve thousand armed for war.
NUM|31|6|And Moses sent them to the war, a thousand from each tribe, together with Phinehas the son of Eleazar the priest, with the vessels of the sanctuary and the trumpets for the alarm in his hand.
NUM|31|7|They warred against Midian, as the LORD commanded Moses, and killed every male.
NUM|31|8|They killed the kings of Midian with the rest of their slain, Evi, Rekem, Zur, Hur, and Reba, the five kings of Midian. And they also killed Balaam the son of Beor with the sword.
NUM|31|9|And the people of Israel took captive the women of Midian and their little ones, and they took as plunder all their cattle, their flocks, and all their goods.
NUM|31|10|All their cities in the places where they lived, and all their encampments, they burned with fire,
NUM|31|11|and took all the spoil and all the plunder, both of man and of beast.
NUM|31|12|Then they brought the captives and the plunder and the spoil to Moses, and to Eleazar the priest, and to the congregation of the people of Israel, at the camp on the plains of Moab by the Jordan at Jericho.
NUM|31|13|Moses and Eleazar the priest and all the chiefs of the congregation went to meet them outside the camp.
NUM|31|14|And Moses was angry with the officers of the army, the commanders of thousands and the commanders of hundreds, who had come from service in the war.
NUM|31|15|Moses said to them, "Have you let all the women live?
NUM|31|16|Behold, these, on Balaam's advice, caused the people of Israel to act treacherously against the LORD in the incident of Peor, and so the plague came among the congregation of the LORD.
NUM|31|17|Now therefore, kill every male among the little ones, and kill every woman who has known man by lying with him.
NUM|31|18|But all the young girls who have not known man by lying with him keep alive for yourselves.
NUM|31|19|Encamp outside the camp seven days. Whoever of you has killed any person and whoever has touched any slain, purify yourselves and your captives on the third day and on the seventh day.
NUM|31|20|You shall purify every garment, every article of skin, all work of goats' hair, and every article of wood."
NUM|31|21|Then Eleazar the priest said to the men in the army who had gone to battle: "This is the statute of the law that the LORD has commanded Moses:
NUM|31|22|only the gold, the silver, the bronze, the iron, the tin, and the lead,
NUM|31|23|everything that can stand the fire, you shall pass through the fire, and it shall be clean. Nevertheless, it shall also be purified with the water for impurity. And whatever cannot stand the fire, you shall pass through the water.
NUM|31|24|You must wash your clothes on the seventh day, and you shall be clean. And afterward you may come into the camp."
NUM|31|25|The LORD said to Moses,
NUM|31|26|"Take the count of the plunder that was taken, both of man and of beast, you and Eleazar the priest and the heads of the fathers' houses of the congregation,
NUM|31|27|and divide the plunder into two parts between the warriors who went out to battle and all the congregation.
NUM|31|28|And levy for the LORD a tribute from the men of war who went out to battle, one out of five hundred, of the people and of the oxen and of the donkeys and of the flocks.
NUM|31|29|Take it from their half and give it to Eleazar the priest as a contribution to the LORD.
NUM|31|30|And from the people of Israel's half you shall take one drawn out of every fifty, of the people, of the oxen, of the donkeys, and of the flocks, of all the cattle, and give them to the Levites who keep guard over the tabernacle of the LORD."
NUM|31|31|And Moses and Eleazar the priest did as the LORD commanded Moses.
NUM|31|32|Now the plunder remaining of the spoil that the army took was 675,000 sheep,
NUM|31|33|72,000 cattle,
NUM|31|34|61,000 donkeys,
NUM|31|35|and 32,000 persons in all, women who had not known man by lying with him.
NUM|31|36|And the half, the portion of those who had gone out in the army, numbered 337,500 sheep,
NUM|31|37|and the LORD's tribute of sheep was 675.
NUM|31|38|The cattle were 36,000, of which the LORD's tribute was 72.
NUM|31|39|The donkeys were 30,500, of which the LORD's tribute was 61.
NUM|31|40|The persons were 16,000, of which the LORD's tribute was 32 persons.
NUM|31|41|And Moses gave the tribute, which was the contribution for the LORD, to Eleazar the priest, as the LORD commanded Moses.
NUM|31|42|From the people of Israel's half, which Moses separated from that of the men who had served in the army-
NUM|31|43|now the congregation's half was 337,500 sheep,
NUM|31|44|36,000 cattle,
NUM|31|45|and 30,500 donkeys,
NUM|31|46|and 16,000 persons-
NUM|31|47|from the people of Israel's half Moses took one of every 50, both of persons and of beasts, and gave them to the Levites who kept guard over the tabernacle of the LORD, as the LORD commanded Moses.
NUM|31|48|Then the officers who were over the thousands of the army, the commanders of thousands and the commanders of hundreds, came near to Moses
NUM|31|49|and said to Moses, "Your servants have counted the men of war who are under our command, and there is not a man missing from us.
NUM|31|50|And we have brought the LORD's offering, what each man found, articles of gold, armlets and bracelets, signet rings, earrings, and beads, to make atonement for ourselves before the LORD."
NUM|31|51|And Moses and Eleazar the priest received from them the gold, all crafted articles.
NUM|31|52|And all the gold of the contribution that they presented to the LORD, from the commanders of thousands and the commanders of hundreds, was 16,750 shekels.
NUM|31|53|(The men in the army had each taken plunder for himself.)
NUM|31|54|And Moses and Eleazar the priest received the gold from the commanders of thousands and of hundreds, and brought it into the tent of meeting, as a memorial for the people of Israel before the LORD.
NUM|32|1|Now the people of Reuben and the people of Gad had a very great number of livestock. And they saw the land of Jazer and the land of Gilead, and behold, the place was a place for livestock.
NUM|32|2|So the people of Gad and the people of Reuben came and said to Moses and to Eleazar the priest and to the chiefs of the congregation,
NUM|32|3|"Ataroth, Dibon, Jazer, Nimrah, Heshbon, Elealeh, Sebam, Nebo, and Beon,
NUM|32|4|the land that the LORD struck down before the congregation of Israel, is a land for livestock, and your servants have livestock."
NUM|32|5|And they said, "If we have found favor in your sight, let this land be given to your servants for a possession. Do not take us across the Jordan."
NUM|32|6|But Moses said to the people of Gad and to the people of Reuben, "Shall your brothers go to the war while you sit here?
NUM|32|7|Why will you discourage the heart of the people of Israel from going over into the land that the LORD has given them?
NUM|32|8|Your fathers did this, when I sent them from Kadesh-barnea to see the land.
NUM|32|9|For when they went up to the Valley of Eshcol and saw the land, they discouraged the heart of the people of Israel from going into the land that the LORD had given them.
NUM|32|10|And the LORD's anger was kindled on that day, and he swore, saying,
NUM|32|11|'Surely none of the men who came up out of Egypt, from twenty years old and upward, shall see the land that I swore to give to Abraham, to Isaac, and to Jacob, because they have not wholly followed me,
NUM|32|12|none except Caleb the son of Jephunneh the Kenizzite and Joshua the son of Nun, for they have wholly followed the LORD.'
NUM|32|13|And the LORD's anger was kindled against Israel, and he made them wander in the wilderness forty years, until all the generation that had done evil in the sight of the LORD was gone.
NUM|32|14|And behold, you have risen in your fathers' place, a brood of sinful men, to increase still more the fierce anger of the LORD against Israel!
NUM|32|15|For if you turn away from following him, he will again abandon them in the wilderness, and you will destroy all this people."
NUM|32|16|Then they came near to him and said, "We will build sheepfolds here for our livestock, and cities for our little ones,
NUM|32|17|but we will take up arms, ready to go before the people of Israel, until we have brought them to their place. And our little ones shall live in the fortified cities because of the inhabitants of the land.
NUM|32|18|We will not return to our homes until each of the people of Israel has gained his inheritance.
NUM|32|19|For we will not inherit with them on the other side of the Jordan and beyond, because our inheritance has come to us on this side of the Jordan to the east."
NUM|32|20|So Moses said to them, "If you will do this, if you will take up arms to go before the LORD for the war,
NUM|32|21|and every armed man of you will pass over the Jordan before the LORD, until he has driven out his enemies from before him
NUM|32|22|and the land is subdued before the LORD; then after that you shall return and be free of obligation to the LORD and to Israel, and this land shall be your possession before the LORD.
NUM|32|23|But if you will not do so, behold, you have sinned against the LORD, and be sure your sin will find you out.
NUM|32|24|Build cities for your little ones and folds for your sheep, and do what you have promised."
NUM|32|25|And the people of Gad and the people of Reuben said to Moses, "Your servants will do as my lord commands.
NUM|32|26|Our little ones, our wives, our livestock, and all our cattle, shall remain there in the cities of Gilead,
NUM|32|27|but your servants will pass over, every man who is armed for war, before the LORD to battle, as my lord orders."
NUM|32|28|So Moses gave command concerning them to Eleazar the priest and to Joshua the son of Nun and to the heads of the fathers' houses of the tribes of the people of Israel.
NUM|32|29|And Moses said to them, "If the people of Gad and the people of Reuben, every man who is armed to battle before the LORD, will pass with you over the Jordan and the land shall be subdued before you, then you shall give them the land of Gilead for a possession.
NUM|32|30|However, if they will not pass over with you armed, they shall have possessions among you in the land of Canaan."
NUM|32|31|And the people of Gad and the people of Reuben answered, "What the LORD has said to your servants, we will do.
NUM|32|32|We will pass over armed before the LORD into the land of Canaan, and the possession of our inheritance shall remain with us beyond the Jordan."
NUM|32|33|And Moses gave to them, to the people of Gad and to the people of Reuben and to the half-tribe of Manasseh the son of Joseph, the kingdom of Sihon king of the Amorites and the kingdom of Og king of Bashan, the land and its cities with their territories, the cities of the land throughout the country.
NUM|32|34|And the people of Gad built Dibon, Ataroth, Aroer,
NUM|32|35|Atroth-shophan, Jazer, Jogbehah,
NUM|32|36|Beth-nimrah and Beth-haran, fortified cities, and folds for sheep.
NUM|32|37|And the people of Reuben built Heshbon, Elealeh, Kiriathaim,
NUM|32|38|Nebo, and Baal-meon (their names were changed), and Sibmah. And they gave other names to the cities that they built.
NUM|32|39|And the sons of Machir the son of Manasseh went to Gilead and captured it, and dispossessed the Amorites who were in it.
NUM|32|40|And Moses gave Gilead to Machir the son of Manasseh, and he settled in it.
NUM|32|41|And Jair the son of Manasseh went and captured their villages, and called them Havvoth-jair.
NUM|32|42|And Nobah went and captured Kenath and its villages, and called it Nobah, after his own name.
NUM|33|1|These are the stages of the people of Israel, when they went out of the land of Egypt by their companies under the leadership of Moses and Aaron.
NUM|33|2|Moses wrote down their starting places, stage by stage, by command of the LORD, and these are their stages according to their starting places.
NUM|33|3|They set out from Rameses in the first month, on the fifteenth day of the first month. On the day after the Passover, the people of Israel went out triumphantly in the sight of all the Egyptians,
NUM|33|4|while the Egyptians were burying all their firstborn, whom the LORD had struck down among them. On their gods also the LORD executed judgments.
NUM|33|5|So the people of Israel set out from Rameses and camped at Succoth.
NUM|33|6|And they set out from Succoth and camped at Etham, which is on the edge of the wilderness.
NUM|33|7|And they set out from Etham and turned back to Pihahiroth, which is east of Baal-zephon, and they camped before Migdol.
NUM|33|8|And they set out from before Hahiroth and passed through the midst of the sea into the wilderness, and they went a three days' journey in the wilderness of Etham and camped at Marah.
NUM|33|9|And they set out from Marah and came to Elim; at Elim there were twelve springs of water and seventy palm trees, and they camped there.
NUM|33|10|And they set out from Elim and camped by the Red Sea.
NUM|33|11|And they set out from the Red Sea and camped in the wilderness of Sin.
NUM|33|12|And they set out from the wilderness of Sin and camped at Dophkah.
NUM|33|13|And they set out from Dophkah and camped at Alush.
NUM|33|14|And they set out from Alush and camped at Rephidim, where there was no water for the people to drink.
NUM|33|15|And they set out from Rephidim and camped in the wilderness of Sinai.
NUM|33|16|And they set out from the wilderness of Sinai and camped at Kibroth-hattaavah.
NUM|33|17|And they set out from Kibroth-hattaavah and camped at Hazeroth.
NUM|33|18|And they set out from Hazeroth and camped at Rithmah.
NUM|33|19|And they set out from Rithmah and camped at Rimmon-perez.
NUM|33|20|And they set out from Rimmon-perez and camped at Libnah.
NUM|33|21|And they set out from Libnah and camped at Rissah.
NUM|33|22|And they set out from Rissah and camped at Kehelathah.
NUM|33|23|And they set out from Kehelathah and camped at Mount Shepher.
NUM|33|24|And they set out from Mount Shepher and camped at Haradah.
NUM|33|25|And they set out from Haradah and camped at Makheloth.
NUM|33|26|And they set out from Makheloth and camped at Tahath.
NUM|33|27|And they set out from Tahath and camped at Terah.
NUM|33|28|And they set out from Terah and camped at Mithkah.
NUM|33|29|And they set out from Mithkah and camped at Hashmonah.
NUM|33|30|And they set out from Hashmonah and camped at Moseroth.
NUM|33|31|And they set out from Moseroth and camped at Bene-jaakan.
NUM|33|32|And they set out from Bene-jaakan and camped at Hor-haggidgad.
NUM|33|33|And they set out from Hor-haggidgad and camped at Jotbathah.
NUM|33|34|And they set out from Jotbathah and camped at Abronah.
NUM|33|35|And they set out from Abronah and camped at Ezion-geber.
NUM|33|36|And they set out from Ezion-geber and camped in the wilderness of Zin (that is, Kadesh).
NUM|33|37|And they set out from Kadesh and camped at Mount Hor, on the edge of the land of Edom.
NUM|33|38|And Aaron the priest went up Mount Hor at the command of the LORD and died there, in the fortieth year after the people of Israel had come out of the land of Egypt, on the first day of the fifth month.
NUM|33|39|And Aaron was 123 years old when he died on Mount Hor.
NUM|33|40|And the Canaanite, the king of Arad, who lived in the Negeb in the land of Canaan, heard of the coming of the people of Israel.
NUM|33|41|And they set out from Mount Hor and camped at Zalmonah.
NUM|33|42|And they set out from Zalmonah and camped at Punon.
NUM|33|43|And they set out from Punon and camped at Oboth.
NUM|33|44|And they set out from Oboth and camped at Iye-abarim, in the territory of Moab.
NUM|33|45|And they set out from Iyim and camped at Dibon-gad.
NUM|33|46|And they set out from Dibon-gad and camped at Almon-diblathaim.
NUM|33|47|And they set out from Almon-diblathaim and camped in the mountains of Abarim, before Nebo.
NUM|33|48|And they set out from the mountains of Abarim and camped in the plains of Moab by the Jordan at Jericho;
NUM|33|49|they camped by the Jordan from Bethjeshimoth as far as Abel-shittim in the plains of Moab.
NUM|33|50|And the LORD spoke to Moses in the plains of Moab by the Jordan at Jericho, saying,
NUM|33|51|"Speak to the people of Israel and say to them, When you pass over the Jordan into the land of Canaan,
NUM|33|52|then you shall drive out all the inhabitants of the land from before you and destroy all their figured stones and destroy all their metal images and demolish all their high places.
NUM|33|53|And you shall take possession of the land and settle in it, for I have given the land to you to possess it.
NUM|33|54|You shall inherit the land by lot according to your clans. To a large tribe you shall give a large inheritance, and to a small tribe you shall give a small inheritance. Wherever the lot falls for anyone, that shall be his. According to the tribes of your fathers you shall inherit.
NUM|33|55|But if you do not drive out the inhabitants of the land from before you, then those of them whom you let remain shall be as barbs in your eyes and thorns in your sides, and they shall trouble you in the land where you dwell.
NUM|33|56|And I will do to you as I thought to do to them."
NUM|34|1|The LORD spoke to Moses, saying,
NUM|34|2|"Command the people of Israel, and say to them, When you enter the land of Canaan (this is the land that shall fall to you for an inheritance, the land of Canaan as defined by its borders),
NUM|34|3|your south side shall be from the wilderness of Zin alongside Edom, and your southern border shall run from the end of the Salt Sea on the east.
NUM|34|4|And your border shall turn south of the ascent of Akrabbim, and cross to Zin, and its limit shall be south of Kadesh-barnea. Then it shall go on to Hazar-addar, and pass along to Azmon.
NUM|34|5|And the border shall turn from Azmon to the Brook of Egypt, and its limit shall be at the sea.
NUM|34|6|"For the western border, you shall have the Great Sea and its coast. This shall be your western border.
NUM|34|7|"This shall be your northern border: from the Great Sea you shall draw a line to Mount Hor.
NUM|34|8|From Mount Hor you shall draw a line to Lebo-hamath, and the limit of the border shall be at Zedad.
NUM|34|9|Then the border shall extend to Ziphron, and its limit shall be at Hazar-enan. This shall be your northern border.
NUM|34|10|"You shall draw a line for your eastern border from Hazar-enan to Shepham.
NUM|34|11|And the border shall go down from Shepham to Riblah on the east side of Ain. And the border shall go down and reach to the shoulder of the Sea of Chinnereth on the east.
NUM|34|12|And the border shall go down to the Jordan, and its limit shall be at the Salt Sea. This shall be your land as defined by its borders all around."
NUM|34|13|Moses commanded the people of Israel, saying, "This is the land that you shall inherit by lot, which the LORD has commanded to give to the nine tribes and to the half-tribe.
NUM|34|14|For the tribe of the people of Reuben by fathers' houses and the tribe of the people of Gad by their fathers' houses have received their inheritance, and also the half-tribe of Manasseh.
NUM|34|15|The two tribes and the half-tribe have received their inheritance beyond the Jordan east of Jericho, toward the sunrise."
NUM|34|16|The LORD spoke to Moses, saying,
NUM|34|17|"These are the names of the men who shall divide the land to you for inheritance: Eleazar the priest and Joshua the son of Nun.
NUM|34|18|You shall take one chief from every tribe to divide the land for inheritance.
NUM|34|19|These are the names of the men: Of the tribe of Judah, Caleb the son of Jephunneh.
NUM|34|20|Of the tribe of the people of Simeon, Shemuel the son of Ammihud.
NUM|34|21|Of the tribe of Benjamin, Elidad the son of Chislon.
NUM|34|22|Of the tribe of the people of Dan a chief, Bukki the son of Jogli.
NUM|34|23|Of the people of Joseph: of the tribe of the people of Manasseh a chief, Hanniel the son of Ephod.
NUM|34|24|And of the tribe of the people of Ephraim a chief, Kemuel the son of Shiphtan.
NUM|34|25|Of the tribe of the people of Zebulun a chief, Elizaphan the son of Parnach.
NUM|34|26|Of the tribe of the people of Issachar a chief, Paltiel the son of Azzan.
NUM|34|27|And of the tribe of the people of Asher a chief, Ahihud the son of Shelomi.
NUM|34|28|Of the tribe of the people of Naphtali a chief, Pedahel the son of Ammihud.
NUM|34|29|These are the men whom the LORD commanded to divide the inheritance for the people of Israel in the land of Canaan."
NUM|35|1|The LORD spoke to Moses in the plains of Moab by the Jordan at Jericho, saying,
NUM|35|2|"Command the people of Israel to give to the Levites some of the inheritance of their possession as cities for them to dwell in. And you shall give to the Levites pasturelands around the cities.
NUM|35|3|The cities shall be theirs to dwell in, and their pasturelands shall be for their cattle and for their livestock and for all their beasts.
NUM|35|4|The pasturelands of the cities, which you shall give to the Levites, shall reach from the wall of the city outward a thousand cubits all around.
NUM|35|5|And you shall measure, outside the city, on the east side two thousand cubits, and on the south side two thousand cubits, and on the west side two thousand cubits, and on the north side two thousand cubits, the city being in the middle. This shall belong to them as pastureland for their cities.
NUM|35|6|The cities that you give to the Levites shall be the six cities of refuge, where you shall permit the manslayer to flee, and in addition to them you shall give forty-two cities.
NUM|35|7|All the cities that you give to the Levites shall be forty-eight, with their pasturelands.
NUM|35|8|And as for the cities that you shall give from the possession of the people of Israel, from the larger tribes you shall take many, and from the smaller tribes you shall take few; each, in proportion to the inheritance that it inherits, shall give of its cities to the Levites."
NUM|35|9|And the LORD spoke to Moses, saying,
NUM|35|10|"Speak to the people of Israel and say to them, When you cross the Jordan into the land of Canaan,
NUM|35|11|then you shall select cities to be cities of refuge for you, that the manslayer who kills any person without intent may flee there.
NUM|35|12|The cities shall be for you a refuge from the avenger, that the manslayer may not die until he stands before the congregation for judgment.
NUM|35|13|And the cities that you give shall be your six cities of refuge.
NUM|35|14|You shall give three cities beyond the Jordan, and three cities in the land of Canaan, to be cities of refuge.
NUM|35|15|These six cities shall be for refuge for the people of Israel, and for the stranger and for the sojourner among them, that anyone who kills any person without intent may flee there.
NUM|35|16|"But if he struck him down with an iron object, so that he died, he is a murderer. The murderer shall be put to death.
NUM|35|17|And if he struck him down with a stone tool that could cause death, and he died, he is a murderer. The murderer shall be put to death.
NUM|35|18|Or if he struck him down with a wooden tool that could cause death, and he died, he is a murderer. The murderer shall be put to death.
NUM|35|19|The avenger of blood shall himself put the murderer to death; when he meets him, he shall put him to death.
NUM|35|20|And if he pushed him out of hatred or hurled something at him, lying in wait, so that he died,
NUM|35|21|or in enmity struck him down with his hand, so that he died, then he who struck the blow shall be put to death. He is a murderer. The avenger of blood shall put the murderer to death when he meets him.
NUM|35|22|"But if he pushed him suddenly without enmity, or hurled anything on him without lying in wait
NUM|35|23|or used a stone that could cause death, and without seeing him dropped it on him, so that he died, though he was not his enemy and did not seek his harm,
NUM|35|24|then the congregation shall judge between the manslayer and the avenger of blood, in accordance with these rules.
NUM|35|25|And the congregation shall rescue the manslayer from the hand of the avenger of blood, and the congregation shall restore him to his city of refuge to which he had fled, and he shall live in it until the death of the high priest who was anointed with the holy oil.
NUM|35|26|But if the manslayer shall at any time go beyond the boundaries of his city of refuge to which he fled,
NUM|35|27|and the avenger of blood finds him outside the boundaries of his city of refuge, and the avenger of blood kills the manslayer, he shall not be guilty of blood.
NUM|35|28|For he must remain in his city of refuge until the death of the high priest, but after the death of the high priest the manslayer may return to the land of his possession.
NUM|35|29|And these things shall be for a statute and rule for you throughout your generations in all your dwelling places.
NUM|35|30|"If anyone kills a person, the murderer shall be put to death on the evidence of witnesses. But no person shall be put to death on the testimony of one witness.
NUM|35|31|Moreover, you shall accept no ransom for the life of a murderer, who is guilty of death, but he shall be put to death.
NUM|35|32|And you shall accept no ransom for him who has fled to his city of refuge, that he may return to dwell in the land before the death of the high priest.
NUM|35|33|You shall not pollute the land in which you live, for blood pollutes the land, and no atonement can be made for the land for the blood that is shed in it, except by the blood of the one who shed it.
NUM|35|34|You shall not defile the land in which you live, in the midst of which I dwell, for I the LORD dwell in the midst of the people of Israel."
NUM|36|1|The heads of the fathers' houses of the clan of the people of Gilead the son of Machir, son of Manasseh, from the clans of the people of Joseph, came near and spoke before Moses and before the chiefs, the heads of the fathers' houses of the people of Israel.
NUM|36|2|They said, "The LORD commanded my lord to give the land for inheritance by lot to the people of Israel, and my lord was commanded by the LORD to give the inheritance of Zelophehad our brother to his daughters.
NUM|36|3|But if they are married to any of the sons of the other tribes of the people of Israel, then their inheritance will be taken from the inheritance of our fathers and added to the inheritance of the tribe into which they marry. So it will be taken away from the lot of our inheritance.
NUM|36|4|And when the jubilee of the people of Israel comes, then their inheritance will be added to the inheritance of the tribe into which they marry, and their inheritance will be taken from the inheritance of the tribe of our fathers."
NUM|36|5|And Moses commanded the people of Israel according to the word of the LORD, saying, "The tribe of the people of Joseph is right.
NUM|36|6|This is what the LORD commands concerning the daughters of Zelophehad, 'Let them marry whom they think best, only they shall marry within the clan of the tribe of their father.
NUM|36|7|The inheritance of the people of Israel shall not be transferred from one tribe to another, for every one of the people of Israel shall hold on to the inheritance of the tribe of his fathers.
NUM|36|8|And every daughter who possesses an inheritance in any tribe of the people of Israel shall be wife to one of the clan of the tribe of her father, so that every one of the people of Israel may possess the inheritance of his fathers.
NUM|36|9|So no inheritance shall be transferred from one tribe to another, for each of the tribes of the people of Israel shall hold on to its own inheritance.'"
NUM|36|10|The daughters of Zelophehad did as the LORD commanded Moses,
NUM|36|11|for Mahlah, Tirzah, Hoglah, Milcah, and Noah, the daughters of Zelophehad, were married to sons of their father's brothers.
NUM|36|12|They were married into the clans of the people of Manasseh the son of Joseph, and their inheritance remained in the tribe of their father's clan.
NUM|36|13|These are the commandments and the rules that the LORD commanded through Moses to the people of Israel in the plains of Moab by the Jordan at Jericho.
