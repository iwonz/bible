ECCL|1|1|Книга Проповідника, сина Давидового, царя в Єрусалимі.
ECCL|1|2|Наймарніша марнота, сказав Проповідник, наймарніша марнота, марнота усе!
ECCL|1|3|Яка користь людині в усім її труді, який вона робить під сонцем?
ECCL|1|4|Покоління відходить, й покоління приходить, а земля віковічно стоїть!
ECCL|1|5|І сонечко сходить, і сонце заходить, і поспішає до місця свого, де сходить воно.
ECCL|1|6|Віє вітер на південь, і на північ вертається, крутиться, крутиться він та й іде, і на круг свій вертається вітер...
ECCL|1|7|Всі потоки до моря пливуть, але море воно не наповнюється: до місця, ізвідки пливуть, ті потоки вони повертаються, щоб знову плисти!
ECCL|1|8|Повні труду всі речі, людина сказати всього не потрапить! Не насититься баченням око, і не наповниться слуханням ухо...
ECCL|1|9|Що було, воно й буде, і що робилося, буде робитись воно, і немає нічого нового під сонцем!...
ECCL|1|10|Буває таке, що про нього говорять: Дивись, це нове! Та воно вже було від віків, що були перед нами!
ECCL|1|11|Нема згадки про перше, а також про наступне, що буде, про них згадки не буде між тими, що будуть потому...
ECCL|1|12|Я, Проповідник, був царем над Ізраїлем в Єрусалимі.
ECCL|1|13|І поклав я на серце своє, щоб шукати й досліджувати мудрістю все, що робилось під небом. Це праця тяжка, яку дав Бог для людських синів, щоб мозолитись нею.
ECCL|1|14|Я бачив усі справи, що чинились під сонцем: й ось усе це марнота та ловлення вітру!...
ECCL|1|15|Покривленого не направиш, а неіснуючого не полічиш!
ECCL|1|16|Говорив я був з серцем своїм та казав: Ось я велику премудрість набув, Найбільшу за всіх, що до мене над Єрусалимом були. І бачило серце моє всяку мудрість і знання.
ECCL|1|17|І поклав я на серце своє, щоб пізнати премудрість, і пізнати безумство й глупоту, і збагнув я, що й це все то ловлення вітру!...
ECCL|1|18|Бо при многості мудрости множиться й клопіт, хто ж пізнання побільшує, той побільшує й біль!...
ECCL|2|1|Сказав був я в серці своєму: Іди но, хай випробую тебе радістю, і придивись до добра, та й воно ось марнота...
ECCL|2|2|На сміх я сказав: Нерозумний, а на радість: Що робить вона?
ECCL|2|3|Задумав я в серці своєму вином оживляти своє тіло, і провадити мудрістю серце своє, і що буду держатись глупоти, аж поки побачу, що ж добре для людських синів, що робили б під небом за короткого часу свого життя.
ECCL|2|4|Поробив я великі діла: поставив для себе доми, задля себе садив виноградники,
ECCL|2|5|запровадив для себе садки та гаї, і понасаджував в них усіляких дерев овочевих.
ECCL|2|6|Наробив я для себе ставів, щоб поливати із них ліс дерев, що виростали.
ECCL|2|7|Набував я для себе рабів та невільниць, були в мене й домівники. А худоби великої та худоби дрібної було в мене більше, ніж у всіх, що в Єрусалимі до мене були!
ECCL|2|8|Назбирав я собі також срібла та золота, і скарбів царів та провінцій, завів я собі співаків та співачок, і всякі приємнощі людських синів, жінок наложниць.
ECCL|2|9|І звеличувавсь я усе більше та більше, над усіх, що в Єрусалимі до мене були, моя мудрість стояла також при мені.
ECCL|2|10|І всього, чого очі мої пожадали, я їм не відмовлював: я не стримував серця свого від жодної втіхи, бо тішилось серце моє від усякого труду мого, і це була частка моя від усякого труду свого!
ECCL|2|11|Та коли я звернувся до всіх своїх чинів, що їх поробили були мої руки, і до труду, що я потрудився був, роблячи, й ось усе це марнота та ловлення вітру, і немає під сонцем нічого корисного!...
ECCL|2|12|І звернувся я, щоб бачити мудрість, і безум, і дурощі. Бо що зробить людина, що прийде вона по царі? Тільки те, що вона вже зробила!
ECCL|2|13|І я побачив, що є перевага у мудрости над глупотою, як є перевага у світла над темрявою:
ECCL|2|14|у мудрого очі його в голові його, а безглуздий у темряві ходить; та теж я пізнав, що доля одна всім їм трапиться!
ECCL|2|15|І промовив я в серці своєму: Коли доля, яка нерозумному трапиться, трапиться також мені, то нащо тоді я мудрішим ставав? І я говорив був у серці своїм, що марнота й оце...
ECCL|2|16|Не лишається пам'яти про мудрого, як і про нерозумного, на вічні віки, в днях наступних зовсім все забудеться, і мудрий вмирає так само, як і нерозумний...
ECCL|2|17|І життя я зненавидів, бо противний мені кожен чин, що під сонцем він чиниться, бо все це марнота та ловлення вітру!...
ECCL|2|18|І зненавидів я ввесь свій труд, що під сонцем трудився я був, бо його позоставлю людині, що буде вона по мені,
ECCL|2|19|а хто знає, чи мудрий той буде чи нерозумний, хто запанує над цілим трудом моїм, над яким я трудився й змудрів був під сонцем? Це марнота також...
ECCL|2|20|І я обернувся чинити, щоб серце моє прийшло в розпач від усього труда, що чинив я під сонцем...
ECCL|2|21|Бо буває людина, що трудиться з мудрістю, зо знанням та із хистом, та все полишає на долю людині, яка не трудилася в тому: Марнота й оце й зло велике!
ECCL|2|22|Та й що має людина зо всього свойого труда та із клопоту серця свого, що під сонцем працює вона?
ECCL|2|23|Бо всі дні її муки, а смуток робота її, і навіть вночі її серце спокою не знає, теж марнота й оце!...
ECCL|2|24|Нема ліпшого земній людині над те, щоб їсти та пити, і щоб душа її бачила добре із труду свого. Та й оце все, я бачив, воно з руки Бога!
ECCL|2|25|Бо хто буде їсти, і хто споживати спроможе без Нього?
ECCL|2|26|Бо людині, що перед лицем Його добра, дає Він премудрість, і пізнання, і радість; а грішникові Він роботу дає, щоб збирати й громадити, щоб пізніше віддати тому, хто добрий перед Божим лицем. Марнота і це все та ловлення вітру!...
ECCL|3|1|Для всього свій час, і година своя кожній справі під небом:
ECCL|3|2|час родитись і час помирати, час садити і час виривати посаджене,
ECCL|3|3|час вбивати і час лікувати, час руйнувати і час будувати,
ECCL|3|4|час плакати й час реготати, час ридати і час танцювати,
ECCL|3|5|час розкидати каміння і час каміння громадити, час обіймати і час ухилятись обіймів,
ECCL|3|6|час шукати і час розгубити, час збирати і час розкидати,
ECCL|3|7|час дерти і час зашивати, час мовчати і час говорити,
ECCL|3|8|час кохати і час ненавидіти, час війні і час миру!
ECCL|3|9|Яка користь трудящому в тім, над чим трудиться він?
ECCL|3|10|Я бачив роботу, що Бог був дав людським синам, щоб трудились над нею,
ECCL|3|11|усе Він прегарним зробив свого часу, і вічність поклав їм у серце, хоч не розуміє людина тих діл, що Бог учинив, від початку та аж до кінця...
ECCL|3|12|Я знаю, немає нічого в них кращого, як тільки радіти й робити добро у своєму житті.
ECCL|3|13|І отож, як котрий чоловік їсть та п'є і в усім своїм труді радіє добром, це дар Божий!
ECCL|3|14|Я знаю, що все, що Бог робить, воно зостається навіки, до того не можна нічого додати, і з того не можна нічого відняти, і Бог так зробив, щоб боялись Його!
ECCL|3|15|Що є, то було вже воно, і що статися має було вже, бо минуле відновлює Бог!
ECCL|3|16|І я бачив під сонцем іще: місце суду, а в нім беззаконня, і місце правди, у ньому ж неправда...
ECCL|3|17|Я сказав був у серці своєму: Судитиме Бог справедливого й несправедливого, бо для кожної справи є час, і на всяке там діло.
ECCL|3|18|Я сказав був у серці своєму: Це для людських синів, щоб Бог випробовував їх, і щоб бачити їм, що вони як ті звірі,
ECCL|3|19|бо доля для людських синів і доля звірини однакова доля для них: як оці помирають, так само вмирають і ті, і для всіх один подих, і нема над твариною вищости людям, марнота бо все!...
ECCL|3|20|Все до місця одного йде: все постало із пороху, і вернеться все знов до пороху...
ECCL|3|21|Хто те знає, чи дух людських синів підіймається вгору, і чи спускається вділ до землі дух скотини?
ECCL|3|22|І я бачив, нема чоловікові кращого, як ділами своїми радіти, бо це доля його! Бо хто поведе його глянути, що буде по ньому?...
ECCL|4|1|І знов я побачив всі утиски, що чинились під сонцем, і сльоза ось утискуваних, та немає для них потішителя, і насилля з руки, що їх гноблять, і немає для них потішителя...
ECCL|4|2|І я похвалив тих померлих, що давно повмирали, більш від живих, що живуть дотепер...
ECCL|4|3|А краще від них від обох тій людині, що досі іще не була, що не бачила чину лихого, що робився під сонцем!
ECCL|4|4|І я бачив ввесь труд та ввесь успіх учинку, викликає заздрість одного до одного, і це все марнота та ловлення вітру!...
ECCL|4|5|Нерозумний сидить, склавши руки свої, та жере своє тіло,
ECCL|4|6|краща повна долоня спокою за повні дві жмені клопоту та за ловлення вітру!...
ECCL|4|7|І знову я бачив марноту під сонцем:
ECCL|4|8|Буває самотній, і не має нікого він іншого, сина чи брата у нього нема, та немає кінця всьому зусиллю його, і не насититься око багатством його, і він не повість: Та для кого дбаю і позбавляю добра свою душу? Марнота й оце, і даремна робота воно...
ECCL|4|9|Краще двом, як одному, бо мають хорошу заплату за труд свій,
ECCL|4|10|і якби вони впали, підійме одне свого друга! Та горе одному, як він упаде, й нема другого, щоб підвести його...
ECCL|4|11|Також коли вдвох покладуться, то тепло їм буде, а як же зогрітись одному?
ECCL|4|12|А коли б хто напав на одного, то вдвох вони стануть на нього, і нитка потрійна не скоро пірветься!
ECCL|4|13|Ліпший убогий та мудрий юнак, аніж цар старий та нерозумний, що вже осторог не приймає,
ECCL|4|14|бо виходить юнак і з в'язниці, щоб зацарювати, хоч у царстві своїм народивсь він убогим!
ECCL|4|15|Я бачив усіх живих, що ходять під сонцем, на боці цього юнака, цього другого, що став він на місце його.
ECCL|4|16|Немає кінця всьому людові, всьому, що був перед ним, та й наступні не втішаться ним, бо й це теж марнота та ловлення вітру!...
ECCL|5|1|(4-17) Пильнуй за ногою своєю, як до Божого дому йдеш, бо прийти, щоб послухати, це краще за жертву безглуздих, бо не знають нічого вони, окрім чинення зла!
ECCL|5|2|(5-1) Не квапся своїми устами, і серце твоє нехай не поспішає казати слова перед Божим лицем, Бог бо на небі, а ти на землі, тому то нехай нечисленними будуть слова твої!
ECCL|5|3|(5-2) Бо як сон наступає через велику роботу, так багато слів має і голос безглуздого.
ECCL|5|4|(5-3) Коли зробиш обітницю Богові, то не зволікай її виповнити, бо в Нього нема уподобання до нерозумних, а що ти обітуєш, сповни!
ECCL|5|5|(5-4) Краще не дати обіту, ніж дати обіт і не сповнити!
ECCL|5|6|(5-5) Не давай своїм устам впроваджувати своє тіло у гріх, і не говори перед Анголом Божим: Це помилка! Пощо Бог буде гніватися на твій голос, і діла твоїх рук буде нищити?
ECCL|5|7|(5-6) Бо марнота в численності снів, як і в многості слів, але ти бійся Бога!
ECCL|5|8|(5-7) Якщо ти побачиш у краї якому утискування бідаря та порушення права та правди, не дивуйся тій речі, бо високий пильнує згори над високим, а над ними Всевишній.
ECCL|5|9|(5-8) І пожиток землі є для всіх, бо поле й сам цар обробляє.
ECCL|5|10|(5-9) Хто срібло кохає, той не насититься сріблом, хто ж кохає багатство з прибутком, це марнота також!
ECCL|5|11|(5-10) Як маєток примножується, то множаться й ті, що його поїдають, і яка користь його власникові, як тільки, щоб бачили очі його?
ECCL|5|12|(5-11) Сон солодкий в трудящого, чи багато, чи мало він їсть, а ситість багатого спати йому не дає.
ECCL|5|13|(5-12) Є лихо болюче, я бачив під сонцем його: багатство, яке бережеться його власникові на лихо йому,
ECCL|5|14|(5-13) і гине багатство таке в нещасливім випадку, а родиться син і немає нічого у нього в руці:
ECCL|5|15|(5-14) як він вийшов нагий із утроби матері своєї, так відходить ізнов, як прийшов, і нічого не винесе він з свого труду, що можна б узяти своєю рукою!...
ECCL|5|16|(5-15) І це теж зло болюче: так само, як він був прийшов, так відійде, і яка йому користь, що трудився на вітер?
ECCL|5|17|(5-16) А до того всі дні свої їв у темноті, і багато мав смутку, й хвороби та люті...
ECCL|5|18|(5-17) Оце, що я бачив, як добре та гарне: щоб їла людина й пила, і щоб бачила добре в усьому своєму труді, що під сонцем ним трудиться в час нечисленних тих днів свого віку, які Бог їй дав, бо це доля її!
ECCL|5|19|(5-18) Також кожна людина, що Бог дав їй багатство й маєтки, і владу їй дав споживати із того, та брати свою частку та тішитися своїм трудом, то це Божий дарунок!
ECCL|5|20|(5-19) Бо вона днів свого життя небагато на пам'яті матиме, то Бог в її серце шле радість!
ECCL|6|1|Є ще зло, що я бачив під сонцем, і багато його між людьми:
ECCL|6|2|Ось людина, що Бог їй багатство дає, і маєтки та славу, і недостатку ні в чому, чого зажадає, не чує вона для своєї душі, але Бог не дав влади їй те споживати, бо чужа людина те поїсть: Це марнота й недуга тяжка!...
ECCL|6|3|Якби сотню дітей наплодив чоловік, і прожив пречисленні літа, і дні віку його були довгі, але не наситилась добрим душа його, а до того не мав би й належного похорону, то кажу: недоноскові краще від нього!...
ECCL|6|4|Бо в марноті прийшов він, і в темряву йде, і в темряві сховане буде імення його,
ECCL|6|5|ані сонця не бачив він, ані пізнав: йому спокійніше від того!...
ECCL|6|6|А коли б він жив двічі по тисячі літ, та не бачив добра, то хіба не до місця одного все йде?
ECCL|6|7|Увесь труд людини для рота її, і пожадання її не виповнюються.
ECCL|6|8|Бо що більшого має мудрець, ніж безглуздий, що має убогий над те, що перед живими уміє ходити?
ECCL|6|9|Краще бачити очима, аніж мандрувати жаданнями, і також це марнота та ловлення вітру...
ECCL|6|10|Що було, тому ймення його вже надане давно, і відоме, що він чоловік, і він не може правуватися з сильнішим від нього,
ECCL|6|11|бо багато речей, що марноту примножуть, але яка користь від них для людини?
ECCL|6|12|Бо хто знає, що добре людині в житті, за небагатьох днів марного життя її, які пробуває вона, немов тінь? Та й що хто розкаже людині, що буде під сонцем по ній?
ECCL|7|1|Краще добре ім'я від оливи хорошої, а день смерти людини від дня її вродження!
ECCL|7|2|Краще ходити до дому жалоби, ніж ходити до дому бенкету, бо то кінець кожній людині, і живий те до серця свого бере!
ECCL|7|3|Кращий смуток від сміху, бо при обличчі сумнім добре серце!
ECCL|7|4|Серце мудрих у домі жалоби, а серце безглуздих у домі веселощів.
ECCL|7|5|Краще слухати докір розумного, аніж слухати пісні безумних,
ECCL|7|6|бо як тріскот тернини під горщиком, такий сміх нерозумного. Теж марнота й оце!...
ECCL|7|7|Коли мудрий кого утискає, то й сам нерозумним стає, а хабар губить серце.
ECCL|7|8|Кінець діла ліпший від початку його; ліпший терпеливий від чванькуватого!
ECCL|7|9|Не спіши в своїм дусі, щоб гніватися, бо гнів спочиває у надрах глупців.
ECCL|7|10|Не кажи: Що це сталось, що перші дні були кращі за ці? бо не з мудрости ти запитався про це.
ECCL|7|11|Добра мудрість з багатством, а прибуток для тих, хто ще сонечко бачить,
ECCL|7|12|бо в тіні мудрости як у тіні срібла, та користь пізнання у тому, що мудрість життя зберігає тому, хто має її.
ECCL|7|13|Розваж Божий учинок, бо хто може те випростати, що Він покривив?
ECCL|7|14|За доброго дня користай із добра, за злого ж розважуй: Одне й друге вчинив Бог на те, щоб людина нічого по собі не знайшла!
ECCL|7|15|В днях марноти своєї я всього набачивсь: буває справедливий, що гине в своїй справедливості, буває й безбожний, що довго живе в своїм злі.
ECCL|7|16|Не будь справедливим занадто, і не роби себе мудрим над міру: пощо нищити маєш себе?
ECCL|7|17|Не будь несправедливим занадто, і немудрим не будь: пощо маєш померти в нечасі своїм?
ECCL|7|18|Добре, щоб ти ухопився за це, але й з того своєї руки не спускай, бо богобоязний втече від усього того.
ECCL|7|19|Мудрість робить мудрого сильнішим за десятьох володарів, що в місті.
ECCL|7|20|Немає людини праведної на землі, що робила б добро й не грішила,
ECCL|7|21|тому не клади свого серця на всякі слова, що говорять, щоб не чути свого раба, коли він лихословить тебе,
ECCL|7|22|знає бо серце твоє, що багато разів також ти лихословив на інших!
ECCL|7|23|Усе це я в мудрості випробував, і сказав: Стану мудрим! Та далека від мене вона!
ECCL|7|24|Далеке оте, що було, і глибоке, глибоке, хто знайде його?
ECCL|7|25|Звернувся я серцем своїм, щоб пізнати й розвідати, та шукати премудрість і розум, та щоб пізнати, що безбожність глупота, а нерозум безумство!
ECCL|7|26|І знайшов я річ гіршу від смерти то жінку, бо пастка вона, її ж серце тенета, а руки її то кайдани!... Хто добрий у Бога врятований буде від неї, а грішного схопить вона!
ECCL|7|27|Подивися, оце я знайшов, сказав Проповідник: рівняймо одне до одного, щоб знайти зрозуміння!
ECCL|7|28|Чого ще шукала душа моя, та не знайшла: я людину знайшов одну з тисячі, але жінки між ними всіма не знайшов!...
ECCL|7|29|Крім того, поглянь, що знайшов я: що праведною вчинив Бог людину, та вигадок усяких шукають вони!...
ECCL|8|1|Хто, як той мудрий, і значення речі хто знає? Розсвітлює мудрість людини обличчя її, і суворість лиця її змінюється.
ECCL|8|2|Я раджу: Наказа царського виконуй, і то ради присяги перед Богом.
ECCL|8|3|Не квапся від нього відходити, не стій при злій справі, бо все, що захоче, він зробить,
ECCL|8|4|бо слово цареве то влада, і хто йому скаже: Що робиш?
ECCL|8|5|Хто виконує заповідь, той не пізнає нічого лихого, серце ж мудрого знає час і право.
ECCL|8|6|Бо для кожної речі час і право своє, бо лихо людини численне на ній,
ECCL|8|7|бо не знає, що буде, і як саме буде, хто їй розповість?
ECCL|8|8|Немає людини, яка панувала б над вітром, щоб стримати вітер, і влади нема над днем смерти, і на війні нема звільнення, і пана свого не врятує безбожність.
ECCL|8|9|Усе це я бачив, і серце своє прикладав я до кожного чину, що відбувався під сонцем. І був час, коли запанувала людина над людиною на лихо для неї.
ECCL|8|10|І я бачив безбожних похованих, і до їхнього гробу приходили, а ті, що чинили добро, повикидані з місця святого, і в місті забуті... Марнота й оце!
ECCL|8|11|Що скоро не чиниться присуд за вчинок лихий, тому серце людських синів повне ними, щоб чинити лихе.
ECCL|8|12|Хоч сто раз чинить грішний лихе, а Бог суд відкладає йому, однако я знаю, що тим буде добре, хто Бога боїться, хто перед обличчям Його має страх!
ECCL|8|13|А безбожному добре не буде, і мов тінь, довгих днів він не матиме, бо він перед Божим лицем страху не має!
ECCL|8|14|Є марнота, яка на землі діється, що є справедливі, що лихо спадає на них, мов за вчинок безбожних, а є безбожні, що добро спадає на них, мов за чин справедливих! Я сказав, що марнота й оце!...
ECCL|8|15|І радість я похваляв: що немає людині під сонцем добра, хіба тільки щоб їсти, та пити та тішитися, і оце супроводить її в її праці за часу життя її, що під сонцем Бог дав був їй.
ECCL|8|16|Коли я поклав своє серце, щоб мудрість пізнати, і побачити чин, що діється він на землі, бо ні вдень ні вночі сну не бачить людина своїми очима,
ECCL|8|17|і коли я побачив усякий чин Бога, тоді я пізнав, що не може людина збагнути чину, під сонцем учиненого! Тому скільки людина не трудиться, щоб дошукатись цього, то не знайде, і коли й мудрий скаже, що знає, не зможе знайти!...
ECCL|9|1|Ото ж бо все це я до серця свого взяв, і бачило серце моє все оце, що праведні й мудрі та їхні учинки у Божій руці, так само любов чи ненависть: Людина не знає нічого, що є перед нею!
ECCL|9|2|Однакове всім випадає: праведному і безбожному, доброму й чистому та нечистому, і тому, хто жертву приносить, і тому, хто жертви не приносить, як доброму, так і грішникові, тому, хто клянеться, як і тому, хто клятви боїться!...
ECCL|9|3|Оце зле у всім, що під сонцем тим діється, що однакове всім випадає, і серце людських синів повне зла, і за життя їхнього безумство в їхньому серці, а по тому до мертвих відходять...
ECCL|9|4|Хто знаходиться поміж живих, той має надію, бо краще собаці живому, ніж левові мертвому!
ECCL|9|5|Бо знають живі, що помруть, а померлі нічого не знають, і заплати немає вже їм, бо забута і пам'ять про них,
ECCL|9|6|і їхнє кохання, і їхня ненависть, та заздрощі їхні загинули вже, і нема вже їм частки навіки ні в чому, що під сонцем тим діється!...
ECCL|9|7|Тож іди, їж із радістю хліб свій, та з серцем веселим вино своє пий, коли Бог уподобав Собі твої вчинки!
ECCL|9|8|Нехай кожного часу одежа твоя буде біла, і нехай на твоїй голові не бракує оливи!
ECCL|9|9|Заживай життя з жінкою, яку ти кохаєш, по всі дні марноти твоєї, що Бог дав для тебе під сонцем на всі дні марноти твоєї, бо оце твоя доля в житті та в твоєму труді, що під сонцем ним трудишся ти!
ECCL|9|10|Все, що всилі чинити рука твоя, теє роби, бо немає в шеолі, куди ти йдеш, ні роботи, ні роздуму, ані знання, ані мудрости!
ECCL|9|11|Знову я бачив під сонцем, що біг не у скорих, і бій не в хоробрих, а хліб не в премудрих, і не в розумних багатство, ні ласка у знавців, а від часу й нагоди залежні вони!
ECCL|9|12|Бо часу свого людина не знає, мов риби, половлені в пагубну сітку, і мов птахи, захоплені в сільце, так хапаються людські сини за час лиха, коли воно нагло спадає на них!...
ECCL|9|13|Також оцю мудрість я бачив під сонцем, і велика для мене здавалась вона:
ECCL|9|14|Було мале місто, і було в ньому мало людей. І раз прийшов цар великий до нього, й його оточив, і побудував проти нього велику облогу.
ECCL|9|15|Але в ньому знайшлася людина убога, та мудра, і вона врятувала те місто своєю премудрістю, та пізніше ніхто не згадав про цю вбогу людину!
ECCL|9|16|І я говорив: Краща мудрість за силу; однако погорджується мудрість бідного, і не слухаються його слів!
ECCL|9|17|Слова мудрих, почуті в спокої, кращі від крику володаря поміж безглуздими.
ECCL|9|18|Мудрість краща від зброї військової, але один грішник погубить багато добра...
ECCL|10|1|Мертві мухи псують та зашумовують оливу мироварника, так трохи глупоти псує мудрість та славу.
ECCL|10|2|Серце мудрого тягне праворуч, а серце безумного ліворуч.
ECCL|10|3|Коли нерозумний і прямою дорогою йде, йому серця бракує, і всім він говорить, що він нерозумний.
ECCL|10|4|Коли гнів володаря стане на тебе, не лишай свого місця, бо лагідність доводить до прощення навіть великих провин.
ECCL|10|5|Є зло, що я бачив під сонцем, мов помилка, що повстає від володаря:
ECCL|10|6|на великих висотах глупота буває поставлена, а багаті сидять у низині!
ECCL|10|7|Я бачив на конях рабів, князі ж пішки ходили, немов ті раби...
ECCL|10|8|Хто яму копає, той в неї впаде, а хто валить мура, того гадина вкусить.
ECCL|10|9|Хто зносить каміння, пораниться ним; хто дрова рубає, загрожений ними.
ECCL|10|10|Як залізо ступіє, й хтось леза не вигострить, той мусить напружити свою силу, та мудрість зарадить йому!
ECCL|10|11|Коли вкусить гадюка перед закляттям, тоді ворожбит не потрібний.
ECCL|10|12|Слова з уст премудрого милість, а губи безумного нищать його:
ECCL|10|13|початок слів його уст глупота, а кінець його уст зле шаленство.
ECCL|10|14|Нерозумний говорить багато, та не знає людина, що буде; а що буде по ньому, хто скаже йому?
ECCL|10|15|Втомляє безумного праця його, бо не знає й дороги до міста.
ECCL|10|16|Горе, краю, тобі, коли цар твій хлопчина, а владики твої спозаранку їдять!
ECCL|10|17|Щасливий ти, краю, коли син шляхетних у тебе царем, а владики твої своєчасно їдять, як ті мужі, а не як п'яниці!
ECCL|10|18|Від лінощів валиться стеля, а з опущення рук тече дах.
ECCL|10|19|Гостину справляють для радощів, і вином веселиться життя, а за срібло все це можна мати.
ECCL|10|20|Навіть у думці своїй не злослов на царя, і в спальні своїй не кляни багача, небесний бо птах віднесе твою мову, а крилатий розкаже про слово твоє...
ECCL|11|1|Хліб свій пускай по воді, бо по багатьох днях знов знайдеш його.
ECCL|11|2|Давай частку на сім чи й на вісім, бо не знаєш, яке буде зло на землі.
ECCL|11|3|Коли переповняться хмари дощем, то виллють на землю його. А коли деревина на південь впаде чи на північ, залишиться на місці, куди деревина впаде.
ECCL|11|4|Хто вважає на вітер, не буде той сіяти, а хто споглядає на хмари, не буде той жати.
ECCL|11|5|Як не відаєш ти, яка то путь вітру, як кості зростають в утробі вагітної, так не відаєш ти чину Бога, що робить усе.
ECCL|11|6|Сій ранком насіння своє, та й під вечір хай не спочиває рука твоя, не знаєш бо ти, котре вийде на краще тобі, оце чи оте, чи обоє однаково добрі.
ECCL|11|7|І світло солодке, і добре очам сонце бачити,
ECCL|11|8|і коли б людина жила й довгі роки, хай за всіх їх вона тішиться, і хай пам'ятає дні темряви, бо їх буде багато, усе, що надійде, марнота!
ECCL|11|9|Тішся, юначе, своїм молодецтвом, а серце твоє нехай буде веселе за днів молодощів твоїх! І ходи ти дорогами серця свого й видінням очей своїх, але знай, що за все це впровадить тебе Бог до суду!
ECCL|11|10|Тому жени смуток від серця свого, і віддаляй зле від тіла твого, бо й дитинство, і рання життєва зоря то марнота!
ECCL|12|1|І пам'ятай в днях юнацтва свого про свого Творця, аж поки не прийдуть злі дні, й не наступлять літа, про які говорити ти будеш: Для мене вони неприємні!
ECCL|12|2|аж поки не стемніє сонце, і світло, і місяць, і зорі, і не вернуться хмари густі за дощем,
ECCL|12|3|у день, коли затремтять ті, хто дім стереже, і зігнуться мужні, і спинять роботу свою млинарі, бо їх стане мало, і потемніють ті, хто в вікно визирає,
ECCL|12|4|і двері подвійні на вулицю замкнені будуть, як зменшиться гуркіт млина, і голос пташини замовкне, і затихнуть всі дочки співучі,
ECCL|12|5|і будуть боятись високого місця, і жахи в дорозі їм будуть, і мигдаль зацвіте, й обтяжіє кобилка, і загине бажання, бо людина відходить до вічного дому свого, а по вулиці будуть ходити довкола голосільники,
ECCL|12|6|аж поки не пірветься срібний шнурок, і не зломиться кругла посудина з золота, і при джерелі не розіб'ється глек, і не зламається коло, й не руне в криницю...
ECCL|12|7|І вернеться порох у землю, як був, а дух вернеться знову до Бога, що дав був його!
ECCL|12|8|Наймарніша марнота, сказав Проповідник, марнота усе!...
ECCL|12|9|Крім того, що Проповідник був мудрий, він навчав ще народ знання. Він важив та досліджував, склав багато приповістей.
ECCL|12|10|Проповідник пильнував знаходити потрібні слова, і вірно писав правдиві слова.
ECCL|12|11|Слова мудрих немов оті леза в ґірлизі, і мов позабивані цвяхи, складачі ж таких слів, вони дані від одного Пастиря.
ECCL|12|12|А понад те, сину мій, будь обережний: складати багато книжок не буде кінця, а багато навчатися мука для тіла!
ECCL|12|13|Підсумок усього почутого: Бога бійся, й чини Його заповіді, бо належить це кожній людині!
ECCL|12|14|Бо Бог приведе кожну справу на суд, і все потаємне, чи добре воно, чи лихе!
