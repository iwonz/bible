ZECH|1|1|大流士 王第二年八月，耶和華的話臨到 易多 的孫子， 比利家 的兒子 撒迦利亞 先知，說：
ZECH|1|2|「耶和華曾向你們祖先大發烈怒。
ZECH|1|3|你要對 以色列 人說，萬軍之耶和華如此說：你們要轉向我，這是萬軍之耶和華說的，我就轉向你們，這是萬軍之耶和華說的。
ZECH|1|4|不要效法你們的祖先。從前的先知呼叫他們說：『萬軍之耶和華如此說，當回轉離開你們的惡道惡行。』他們卻不聽，也不順從我。這是耶和華說的。
ZECH|1|5|你們的祖先在哪裏呢？那些先知能永遠存活嗎？
ZECH|1|6|然而我的言語和律例，就是我所吩咐我僕人眾先知的，豈不臨到你們的祖先嗎？他們就回轉，說：萬軍之耶和華定意按我們的所作所為對待我們，他也已經照樣行了。」
ZECH|1|7|大流士 第二年十一月，就是細罷特月二十四日，耶和華的話臨到 易多 的孫子， 比利家 的兒子 撒迦利亞 先知，說：
ZECH|1|8|「我夜間觀看，看哪，有一人騎著紅馬，站在窪地的番石榴樹中間。在他身後有紅色、褐色和白色的馬。」
ZECH|1|9|我說：「主啊，這是甚麼意思？」與我說話的天使說：「我要指示你這是甚麼意思。」
ZECH|1|10|那站在番石榴樹中間的人回答說：「這是奉耶和華差遣，在遍地巡邏的。」
ZECH|1|11|他們對站在番石榴樹中間耶和華的使者說：「我們在遍地巡邏，看哪，全地都安息平靜。」
ZECH|1|12|於是，耶和華的使者說：「萬軍之耶和華啊，你惱恨 耶路撒冷 和 猶大 的城鎮已經七十年了，你不施憐憫要到幾時呢？」
ZECH|1|13|耶和華就用美善的話和安慰的話回答那與我說話的天使。
ZECH|1|14|與我說話的天使對我說：「你要宣告，萬軍之耶和華如此說：我為 耶路撒冷 而妒忌，為 錫安 大大妒忌。
ZECH|1|15|我非常惱怒那享安逸的列國，因我從前稍微惱怒，他們就越發加害。
ZECH|1|16|所以耶和華如此說：現在我回到 耶路撒冷 ，仍要施憐憫，我的殿要重建在其中，準繩必拉在 耶路撒冷 之上。這是萬軍之耶和華說的。
ZECH|1|17|你要再宣告，萬軍之耶和華如此說：我的城鎮要再度繁榮發達。耶和華必再安慰 錫安 ，揀選 耶路撒冷 。」
ZECH|1|18|我舉目觀看，看哪，有四隻角。
ZECH|1|19|我問那與我說話的天使：「這是甚麼意思？」他對我說：「這是擊散 猶大 、 以色列 和 耶路撒冷 的角。」
ZECH|1|20|耶和華又把四個匠人指給我看。
ZECH|1|21|我問：「這些人來做甚麼呢？」他說：「那是擊散 猶大 的角，使人不敢抬頭；但這些匠人前來威嚇列國，打掉列國的角，因為他們舉起角來擊散 猶大 地。」
ZECH|2|1|我舉目觀看，看哪，有一人手拿丈量的繩。
ZECH|2|2|我問：「你到哪裏去？」他對我說：「要去丈量 耶路撒冷 ，看有多寬多長。」
ZECH|2|3|看哪，與我說話的天使出去 ，另有一位天使迎著他來，
ZECH|2|4|對他說：「你跑去告訴這個年輕人說， 耶路撒冷 必有人居住，如同無城牆的鄉村，因為其中的人和牲畜很多。
ZECH|2|5|耶和華說：『我要作 耶路撒冷 四圍火的城牆，並要作城中的榮耀。』」
ZECH|2|6|耶和華說：「來，來！你們要從北方之地逃回；因我曾把你們分散到天的四方 。這是耶和華說的。」
ZECH|2|7|來！住 巴比倫 的 錫安 百姓啊，逃吧！
ZECH|2|8|萬軍之耶和華在顯出榮耀之後，差遣我到擄掠你們的列國那裏，他如此說：「碰你們的就是碰他自己 眼中的瞳人。
ZECH|2|9|看哪，我要揮手攻擊他們，他們就必作自己奴僕的擄物。」你們就知道萬軍之耶和華差遣了我。
ZECH|2|10|耶和華說：「 錫安 哪，應當歡樂歌唱，因為，看哪，我要來，要住在你中間。
ZECH|2|11|在那日，必有許多國家歸附耶和華，作我的子民。我要住 在你中間。」你就知道萬軍之耶和華差遣我到你那裏去。
ZECH|2|12|耶和華必收回 猶大 ，作為他聖地的產業，他必再度揀選 耶路撒冷 。
ZECH|2|13|凡血肉之軀都當在耶和華面前靜默無聲，因為他從他的聖所奮起了。
ZECH|3|1|天使 指給我看： 約書亞 大祭司站在耶和華的使者面前，撒但站在 約書亞 的右邊控告他。
ZECH|3|2|耶和華向撒但說：「撒但哪，耶和華責備你！揀選 耶路撒冷 的耶和華責備你！這不是從火中抽出來的一根柴嗎？」
ZECH|3|3|約書亞 穿著污穢的衣服，站在那使者面前。
ZECH|3|4|使者吩咐那些侍立在他面前的說：「脫去他污穢的衣服。」又對 約書亞 說：「你看，我使你的罪孽離開你，要給你穿上華美的衣服。」
ZECH|3|5|我說 ：「要將潔淨的冠冕戴在他頭上。」他們就把潔淨的冠冕戴在他頭上，給他穿上華美的衣服，耶和華的使者在旁邊站立。
ZECH|3|6|耶和華的使者告誡 約書亞 說，
ZECH|3|7|萬軍之耶和華如此說：「你若遵行我的道，謹守我的命令，就可以管理我的家，看守我的院宇；我也要使你在這些侍立的人中間來往。
ZECH|3|8|約書亞 大祭司啊，你和坐在你面前的同伴都當聽，因為他們是作預兆的：看哪，我必使我僕人 大衛 的苗裔 長出。
ZECH|3|9|看哪，這是我在 約書亞 面前所立的石頭，這一塊石頭上有七眼。看哪，我要親自雕刻這石頭，並在一日之間除掉這地的罪孽。這是萬軍之耶和華說的。
ZECH|3|10|在那日，你們各人要請鄰舍坐在葡萄樹和無花果樹下。這是萬軍之耶和華說的。」
ZECH|4|1|那與我說話的天使又來叫醒我，好像人睡覺時被喚醒一樣。
ZECH|4|2|他問我：「你看見甚麼？」我說：「我看見了，看哪，有一個純金的燈臺，頂上有燈座，其上有七盞燈，每盞燈的上頭有七根管子；
ZECH|4|3|旁邊有兩棵橄欖樹，一棵在燈座的右邊，一棵在燈座的左邊。」
ZECH|4|4|我問與我說話的天使說：「主啊，這是甚麼意思？」
ZECH|4|5|與我說話的天使回答，對我說：「你不知道這是甚麼意思嗎？」我說：「主啊，我不知道。」
ZECH|4|6|他回答我說：「這是耶和華指示 所羅巴伯 的話。萬軍之耶和華說：不是倚靠勢力，不是倚靠才能，乃是倚靠我的靈方能成事 。
ZECH|4|7|大山哪，你算甚麼呢？在 所羅巴伯 面前，你必夷為平地。他安放頂上的那塊石頭，人就歡呼：『願恩惠、恩惠歸與這殿！』」
ZECH|4|8|耶和華的話臨到我，說：
ZECH|4|9|「 所羅巴伯 的手立了這殿的根基，他的手也必完成這工，你就知道萬軍之耶和華差遣我到你們這裏。
ZECH|4|10|誰藐視這日的事為小呢？他們見 所羅巴伯 手拿石垂線就歡喜。這七盞燈 是耶和華的眼睛，遍察全地。」
ZECH|4|11|我問天使說：「那麼在燈臺左右的這兩棵橄欖樹是甚麼意思呢？」
ZECH|4|12|我再次問他：「這兩根橄欖樹枝在兩根流出金色油的金嘴旁邊，是甚麼意思呢？」
ZECH|4|13|他對我說：「你不知道這是甚麼意思嗎？」我說：「主啊，我不知道。」
ZECH|4|14|他說：「這是兩位受膏者，侍立在全地之主的旁邊。」
ZECH|5|1|我又舉目觀看，看哪，有一飛行的書卷。
ZECH|5|2|他問我：「你看見甚麼？」我回答：「我看見一飛行的書卷，長二十肘，寬十肘。」
ZECH|5|3|他對我說：「這就是向全地面發出的詛咒。凡偷竊的必按書卷這面的話除滅，凡起假誓的必按書卷那面的話除滅。
ZECH|5|4|萬軍之耶和華說：我要把這書卷送出去，進入偷竊者的家和指著我名起假誓者的家，停留在他家裏，連房屋帶木頭和石頭都毀滅了。」
ZECH|5|5|與我說話的天使前來，對我說：「你要舉目觀看，看那出現的是甚麼。」
ZECH|5|6|我問：「這是甚麼呢？」他說：「這出現的是量器 。」又說：「是他們的眼目，遍行全地 。」
ZECH|5|7|看哪，圓形的鉛蓋被抬起來，有一個婦人坐在量器中。
ZECH|5|8|天使說：「這是罪惡。」他就把婦人推進量器裏，把鉛蓋壓在量器的口上。
ZECH|5|9|於是我舉目觀看，看哪，有兩個婦人前來，她們的翅膀中有風，翅膀如同鸛鳥的翅膀。她們把量器抬起來，懸在天地之間。
ZECH|5|10|我問那與我說話的天使：「她們要把量器抬到哪裏去呢？」
ZECH|5|11|他對我說：「要抬到 示拿 地去，為它建造房屋；等預備妥當，就把它安放在自己的臺座上。」
ZECH|6|1|我又舉目觀看，看哪，有四輛馬車從兩座山的中間出來；那兩座山是銅山。
ZECH|6|2|第一輛車套著紅馬，第二輛車套著黑馬，
ZECH|6|3|第三輛車套著白馬，第四輛車套著帶斑點的馬，都是強壯的 。
ZECH|6|4|我就回應與我說話的天使說：「主啊，這是甚麼意思？」
ZECH|6|5|天使回答，對我說：「這是天的四風，是從全地之主面前出來的。」
ZECH|6|6|套著黑馬的車往北方之地去，白馬跟隨在後；有斑點的馬往南方之地去；
ZECH|6|7|那些壯馬出來，急著要在地上巡邏。天使說：「你們只管在地上巡邏。」牠們就在地上巡邏。
ZECH|6|8|他又呼叫我，告訴我說：「你看，往北方地去的已在北方之地使我放心。」
ZECH|6|9|耶和華的話臨到我，說：
ZECH|6|10|「你要拿從 巴比倫 歸來的被擄之人 黑玳 、 多比雅 、 耶大雅 所獻的，當日就要進到 西番雅 的兒子 約西亞 的家裏，
ZECH|6|11|拿這金銀做冠冕，戴在 約撒答 的兒子 約書亞 大祭司的頭上；
ZECH|6|12|對他說，萬軍之耶和華如此說：『看哪，那名稱為 大衛 苗裔的，要在本處生長，並要建造耶和華的殿。
ZECH|6|13|就是他，要建造耶和華的殿，他要承受尊榮，坐在位上掌王權；又有一位祭司坐在自己的位上，兩職之間籌劃和平。
ZECH|6|14|這冠冕要歸 希連 、 多比雅 、 耶大雅 ，和 西番雅 的兒子 賢 ，放在耶和華的殿裏作為紀念。』」
ZECH|6|15|遠方的人要來建造耶和華的殿，你們因此就知道，萬軍之耶和華差遣我到你們這裏來。你們若留意聽從耶和華－你們上帝的話，這事必然成就。
ZECH|7|1|大流士 王第四年九月，就是基斯流月初四，耶和華的話臨到 撒迦利亞 。
ZECH|7|2|那時 伯特利 人已經差遣 沙利色 和 利堅‧米勒 ，並他們的人，去懇求耶和華的恩，
ZECH|7|3|問萬軍之耶和華殿中的祭司，又問先知：「我當如歷年以來所行，在五月哭泣齋戒嗎？」
ZECH|7|4|萬軍之耶和華的話臨到我，說：
ZECH|7|5|「你要向這地全體百姓和祭司說：『你們這七十年來，在五月、七月禁食悲哀，豈是真的向我禁食嗎？
ZECH|7|6|你們吃喝，不是為自己吃，為自己喝嗎？
ZECH|7|7|當 耶路撒冷 和四圍的城鎮有人居住，享繁榮， 尼革夫 和 謝非拉 也有人居住的時候，耶和華藉從前的先知所宣告的，你們不當聽嗎？』」
ZECH|7|8|耶和華的話臨到 撒迦利亞 ，說：
ZECH|7|9|「萬軍之耶和華如此說：你們要按真正的公平來審判，彼此以慈愛憐憫相待。
ZECH|7|10|不可欺壓寡婦、孤兒、寄居的和困苦的人。誰都不可心裏謀害弟兄。
ZECH|7|11|他們卻不留意；聳肩悖逆，耳朵發沉，不肯聽從。
ZECH|7|12|他們的心堅硬如金剛石，不聽律法和萬軍之耶和華藉著他的靈差遣從前先知所說的話。因此，萬軍之耶和華大發烈怒。
ZECH|7|13|萬軍之耶和華說：我曾呼喚他們，他們不聽；將來他們呼求我，我也不聽！
ZECH|7|14|我必以旋風將他們吹散到素不認識的萬國中。他們離開以後，地就荒涼，無人來往經過；他們使美好之地荒涼了。」
ZECH|8|1|萬軍之耶和華的話臨到我，說：
ZECH|8|2|「萬軍之耶和華如此說：我為 錫安 而妒忌，大大妒忌；我為了它妒忌而大發烈怒。
ZECH|8|3|耶和華如此說：我要回到 錫安 ，住在 耶路撒冷 中間。 耶路撒冷 必稱為忠實的城，萬軍之耶和華的山必稱為聖山。
ZECH|8|4|萬軍之耶和華如此說：將來必有年老的男女坐在 耶路撒冷 的廣場上，各人因年紀老邁而手拿枴杖。
ZECH|8|5|城裏的廣場滿有男孩女孩在玩耍。
ZECH|8|6|萬軍之耶和華如此說：在那些日子，即使這事在這餘民眼中看為奇妙，難道在我眼中也看為奇妙嗎？這是萬軍之耶和華說的。
ZECH|8|7|萬軍之耶和華如此說：看哪，我要從日出之地、從日落之地拯救我的子民。
ZECH|8|8|我要領他們來，使他們住在 耶路撒冷 中間。他們要作我的子民，我要作他們的上帝，都憑信實和公義。
ZECH|8|9|「萬軍之耶和華如此說：你們的手要堅強；這些日子，你們已聽見先知的口，在萬軍之耶和華殿的根基立定、聖殿建造的日子所說的這些話。
ZECH|8|10|那些日子以前，人得不著工價，牲畜也無人雇用；且因敵人的緣故，出入不得平安；因我使人與人互相攻擊。
ZECH|8|11|但如今，我對這餘民必不像先前的日子。這是萬軍之耶和華說的。
ZECH|8|12|因為他們要平安撒種，葡萄樹要結果子，土地必有出產，天也必降甘露。我要使這餘民享受這一切。
ZECH|8|13|猶大 家和 以色列 家啊，你們從前在列國中怎樣成為可詛咒的；照樣，我要拯救你們，使你們得福 。不要懼怕，你們的手要堅強。
ZECH|8|14|「萬軍之耶和華如此說：你們祖先惹我發怒的時候，我怎樣定意降禍，並不改變；萬軍之耶和華說，
ZECH|8|15|這些日子我也定意施恩給 耶路撒冷 和 猶大 家；你們不要懼怕。
ZECH|8|16|你們所當行的是這樣：每個人要與鄰舍說誠實話，在城門口要按真正的公平來審判，使人和睦。
ZECH|8|17|誰都不可心裏謀害鄰舍，也不可喜愛起假誓，因為這些事都為我所恨惡。這是耶和華說的。」
ZECH|8|18|萬軍之耶和華的話臨到我，說：
ZECH|8|19|「萬軍之耶和華如此說：四月的禁食、五月的禁食、七月的禁食和十月的禁食，必成為 猶大 家的歡喜和快樂，以及美好的節期；所以你們要喜愛誠實與和平。
ZECH|8|20|「萬軍之耶和華如此說：將來還有眾百姓和許多城鎮的居民要來。
ZECH|8|21|這城的居民必到那城，說：『我們快去懇求耶和華的恩，尋求萬軍之耶和華；我自己也要去。』
ZECH|8|22|必有許多民族和強盛的國家來到 耶路撒冷 尋求萬軍之耶和華，懇求耶和華的恩。
ZECH|8|23|萬軍之耶和華如此說：在那些日子，列國中說各種語言的人，必有十個人強拉住一個 猶大 人衣服的邊，說：『我們要與你們同去，因為我們聽見上帝與你們同在了。』」
ZECH|9|1|耶和華的默示， 他的話臨到 哈得拉 地、 大馬士革 －因世人和 以色列 各支派的眼目都向著耶和華－
ZECH|9|2|和鄰近的 哈馬 ， 以及 推羅 和 西頓 。 因為它極有智慧，
ZECH|9|3|推羅 為自己建造堅固城 ， 堆起銀子如塵沙， 純金如街上的泥土。
ZECH|9|4|看哪，主必趕出它， 重創它海上的勢力， 它必被火吞滅。
ZECH|9|5|亞實基倫 看見必懼怕， 迦薩 看見甚痛苦， 以革倫 因失了盼望而蒙羞； 迦薩 必不再有君王， 亞實基倫 也不再有人居住，
ZECH|9|6|混血的人要住在 亞實突 ； 我必除滅 非利士 人的驕傲。
ZECH|9|7|我要除去他口中帶血之肉 和牙齒內可憎之物。 他必作餘民歸於我們的上帝， 在 猶大 像族長一樣； 以革倫 必如 耶布斯 人。
ZECH|9|8|我要紮營在我的家， 敵軍不得任意往來， 暴虐的人也不再經過， 因為我親眼看顧。
ZECH|9|9|錫安 哪，應當大大喜樂； 耶路撒冷 啊，應當歡呼。 看哪，你的王來到你這裏！ 他是公義的，並且施行拯救， 謙和地騎著驢， 騎著小驢，驢的駒子。
ZECH|9|10|我必除滅 以法蓮 的戰車 和 耶路撒冷 的戰馬； 戰爭的弓也必剪除。 他要向列國講和平； 他的權柄必從這海管到那海， 從 大河 管到地極。
ZECH|9|11|錫安 哪，我因與你立約的血， 要從無水坑裏釋放你中間被囚的人。
ZECH|9|12|被囚而有指望的人哪，要轉回堡壘； 我今日宣告，我必加倍補償你。
ZECH|9|13|我為自己把 猶大 彎緊， 我使 以法蓮 如滿弓。 錫安 哪，我要喚起你的兒女， 希臘 啊，我要攻擊你的兒女， 使你如勇士的刀。
ZECH|9|14|耶和華要顯現在他們身上， 他的箭要射出如閃電。 主耶和華必吹角， 乘南方的旋風而行。
ZECH|9|15|萬軍之耶和華必保護他們； 他們要吞滅，要踐踏彈弓的石頭 ； 他們吶喊，狂飲 如喝酒， 如盛滿的碗， 又如壇的四角。
ZECH|9|16|當那日，耶和華－他們的上帝 必看他的百姓如羊群，拯救他們； 因為他們如冠冕上的寶石， 在他的地上如旗幟高舉 。
ZECH|9|17|他是何等善！ 他是何其美！ 五穀使少男強壯， 新酒使少女健美。
ZECH|10|1|春雨的季節，你們要向耶和華求雨。 耶和華發出雷電， 為眾人降下大雨， 把田園的菜蔬賜給人。
ZECH|10|2|因為家中神像所言的是虛空， 占卜者所見的是虛假， 他們講說假夢， 徒然安慰人。 所以眾人如羊流離， 因無牧人就受欺壓。
ZECH|10|3|我的怒氣向牧人發作， 我必懲罰那為首的 ； 萬軍之耶和華眷顧他的羊群， 就是 猶大 家， 必使他們如戰場上的駿馬。
ZECH|10|4|房角石從他而出， 橛子從他而出， 戰爭的弓也從他而出， 每一個掌權的都從他而出。
ZECH|10|5|他們必如戰場上的勇士， 踐踏仇敵如街上的泥土。 他們必爭戰，因為耶和華與他們同在， 他們必使騎馬的羞愧。
ZECH|10|6|我要堅固 猶大 家， 拯救 約瑟 家， 我要領他們歸回，因我憐憫他們， 他們必像我未曾棄絕他們一樣； 都因我是耶和華－他們的上帝， 我必應允他們。
ZECH|10|7|以法蓮 人必如勇士， 他們心中暢快如同喝酒； 他們的兒女看見就歡喜， 他們的心必因耶和華喜樂。
ZECH|10|8|我要呼叫，聚集他們， 因我已經救贖他們。 他們的人數必增添， 如從前增添一樣。
ZECH|10|9|我要將他們分散在列國中， 他們必在遠方記得我； 他們與兒女都必存活， 他們要歸回。
ZECH|10|10|我必使他們從 埃及 地歸回， 從 亞述 召集他們， 領他們到 基列 地和 黎巴嫩 ； 這些還不夠他們居住。
ZECH|10|11|耶和華 必經過苦海，擊打海浪。 尼羅河 的深處全都枯乾， 亞述 的驕傲必降卑， 埃及 的權杖必除去。
ZECH|10|12|我要使他們倚靠耶和華，得以堅固， 他們必奉他的名而行 ； 這是耶和華說的。
ZECH|11|1|黎巴嫩 哪，敞開你的門， 任火吞滅你的香柏樹。
ZECH|11|2|哀號吧，松樹！ 因為香柏樹傾倒了，高大的樹毀壞了。 哀號吧， 巴珊 的橡樹！ 因為茂盛的樹林倒下來了。
ZECH|11|3|聽啊，有牧人在哀號， 因他們的榮華敗落了； 聽啊，有少壯獅子咆哮， 因 約旦河 旁的叢林荒廢了。
ZECH|11|4|耶和華－我的上帝如此說：「你要牧養這群將宰的羊。
ZECH|11|5|買羊的宰了他們，卻不認為自己有罪；賣他們的也說：『耶和華是應當稱頌的，因我富足了。』牧養他們的並不憐憫他們。
ZECH|11|6|我不再憐憫這地的居民。看哪，我要將這些人交在各人的鄰舍和君王手中；他們必毀滅這地，我卻不救任何一個脫離他們的手。這是耶和華說的。」
ZECH|11|7|於是，我牧養這群將宰的羊，就是羊群中最困苦的 ；我拿著兩根杖，一根我稱為「恩惠」 ，一根稱為「聯合」。這樣，我就牧養這群羊。
ZECH|11|8|一個月之內，我廢除了三個牧人，因為我的心厭煩他們，他們的心也憎惡我。
ZECH|11|9|我就說：「我不牧養你們。要死的，由他死；滅亡的，由他滅亡；剩餘的，由他們彼此吞食。」
ZECH|11|10|我拿起那根稱為「恩惠」的杖，折斷它，表明我廢棄與萬民所立的約。
ZECH|11|11|當日約就廢了。因此，那些羊群中最困苦的 ，看著我，就知道這真是耶和華的話。
ZECH|11|12|我對他們說：「你們若看為美，就給我工價。不然，就罷了！」於是他們秤了三十塊銀錢作為我的工價。
ZECH|11|13|耶和華對我說：「把它丟給窯戶。那是他們對我所估定的好價錢！」我就取這三十塊銀錢，在耶和華的殿中將它丟給窯戶。
ZECH|11|14|我又折斷第二根杖，就是稱為「聯合」的那根杖，表明我廢棄 猶大 與 以色列 弟兄間的情誼。
ZECH|11|15|耶和華對我說：「你再把愚昧牧人所用的器具拿來，
ZECH|11|16|因為，看哪，我要在這地立一個牧人；他不看顧將亡的，不尋找分散的，不醫治受傷的，也不牧養強壯的；卻要吞吃肥羊的肉，撕裂牠們的蹄。
ZECH|11|17|禍哉！無用的牧人丟棄羊群， 刀必臨到他的膀臂和右眼上； 他的膀臂必全然枯乾， 他的右眼也必昏暗失明。」
ZECH|12|1|耶和華的默示，他的話論到 以色列 。 鋪張諸天、建立地基、造人裏面之靈的耶和華說：
ZECH|12|2|「看哪，我要使 耶路撒冷 成為令四圍列國百姓昏醉的杯； 耶路撒冷 被圍困， 猶大 也一樣受困 。
ZECH|12|3|在那日，我要使 耶路撒冷 成為萬民的一塊沉重石頭，凡舉起它的必受重傷；地上的萬國都聚集攻擊它。
ZECH|12|4|到那日，我必令一切的馬匹驚惶，使騎馬的癲狂。我必張開眼睛看顧 猶大 家，卻使列國一切的馬匹瞎眼。這是耶和華說的。
ZECH|12|5|猶大 的族長心裏要說：『 耶路撒冷 的居民因倚靠萬軍之耶和華－他們的上帝，就成為我的力量 。』
ZECH|12|6|「那日，我必使 猶大 的族長如柴堆中的火盆，又如禾捆裏的火把；他們必左右吞滅四圍列國的百姓。 耶路撒冷 卻仍屹立在本處，仍在 耶路撒冷 ！
ZECH|12|7|「耶和華要先拯救 猶大 的帳棚，免得 大衛 家的榮耀和 耶路撒冷 居民的榮耀勝過 猶大 。
ZECH|12|8|那日，耶和華必保護 耶路撒冷 的居民。他們中間軟弱的在那日必如 大衛 ； 大衛 家必如上帝，如行在他們前面的耶和華的使者。
ZECH|12|9|那日，我必定意滅絕前來攻擊 耶路撒冷 的萬國。」
ZECH|12|10|「我要將那施恩與懇求的靈，澆灌 大衛 家和 耶路撒冷 的居民。他們必仰望我，就是他們所扎的那位。他們必為他悲傷，如喪獨子，又為他哀哭，如喪長子。
ZECH|12|11|那日，在 耶路撒冷 必有大大的哀號，如 米吉多 平原上 哈達‧臨門 的哀號。
ZECH|12|12|這地必哀哭：一家一家地哭， 大衛 家的家族聚在一處，他們的婦女聚在一處； 拿單 家的家族聚在一處，他們的婦女聚在一處。
ZECH|12|13|利未 家的家族聚在一處，他們的婦女聚在一處； 示每 家的家族聚在一處，他們的婦女聚在一處。
ZECH|12|14|其餘的各家，每一家的家族聚在一處，他們的婦女聚在一處。」
ZECH|13|1|「在那日，因罪惡與污穢的緣故，必有一泉源為 大衛 家和 耶路撒冷 的居民而開。」
ZECH|13|2|萬軍之耶和華說：「在那日，我要從地上除滅偶像的名，使它不再被記得；我也必使這地不再有先知，不再有污穢的靈。
ZECH|13|3|若還有人說預言，生他的父母必對他說：『你不得存活，因為你假借耶和華的名說謊話。』生他的父母在他說預言時，要將他刺死。
ZECH|13|4|那日，凡作先知說預言的必因所論的異象羞愧，不再穿毛皮外袍哄騙人。
ZECH|13|5|他要說：『我不是先知，我是耕地的；我從幼年就作人的奴僕。』
ZECH|13|6|有人對他說：『你兩手臂間是甚麼傷呢？』他說：『這是我在親友家中所受的傷。』」
ZECH|13|7|萬軍之耶和華說： 刀劍哪，興起攻擊我的牧人， 攻擊我的同伴吧！ 要擊打牧人，羊就分散了； 我必反手攻擊那微小的。
ZECH|13|8|這全地的人， 三分之二將被剪除而死， 三分之一仍必存留。 這是耶和華說的。
ZECH|13|9|我要使這三分之一經過火， 熬煉他們，如熬煉銀子； 試煉他們，如試煉金子。 他們要求告我的名， 我必應允他們。 我說：「這是我的子民。」 他們要說：「耶和華是我的上帝。」
ZECH|14|1|看哪，耶和華的日子臨近了，你的財物必被搶掠，在你中間被瓜分。
ZECH|14|2|我要招聚萬國與 耶路撒冷 爭戰；城必被攻取，房屋被搶奪，婦女被玷污，城中的一半被擄去；但其餘的百姓不會從城中被剪除。
ZECH|14|3|那時，耶和華要出去與那些國家打仗，如同從前戰爭的日子打仗一樣。
ZECH|14|4|那日，他的腳必站在 橄欖山 上，這山面向 耶路撒冷 的東邊。 橄欖山 必從中間裂開，自東至西成為極大的谷；山的一半向北挪移，一半向南挪移。
ZECH|14|5|你們要從我的山谷中逃跑，因為山谷必延到 亞薩 。你們要逃跑，如在 猶大 王 烏西雅 年間逃避大地震一樣 。耶和華－我的上帝必降臨，所有的聖者與你 同來。
ZECH|14|6|在那日，必沒有光，不會放晴，只有烏雲 。
ZECH|14|7|耶和華所知道的那一日，沒有白天，沒有黑夜，到了晚上仍有亮光。
ZECH|14|8|在那日，必有活水從 耶路撒冷 出來，一半往東海流，一半往西海流；冬夏都是如此。
ZECH|14|9|耶和華要作全地的王。那日，耶和華必為獨一無二，他的名也是獨一無二。
ZECH|14|10|從 迦巴 直到 耶路撒冷 南方的 臨門 ，全地要變為曠野。 耶路撒冷 要矗立於本處，從 便雅憫門 到 舊門 ，又到 角門 ，並從 哈楠業樓 ，直到王的酒池。
ZECH|14|11|人要住在其中，不再有詛咒； 耶路撒冷 必安然屹立。
ZECH|14|12|這是耶和華所降的災殃，要攻擊那些與 耶路撒冷 作戰的萬民；他們兩腳站立時，肉要潰爛，眼在眶中潰爛，舌在口中也潰爛。
ZECH|14|13|那日，耶和華必使他們大大混亂。他們彼此用手揪住，用手互相攻擊。
ZECH|14|14|猶大 也要在 耶路撒冷 打仗 。那時四圍各國的財物，就是許許多多的金銀和衣服，必被收聚。
ZECH|14|15|馬匹、騾子、駱駝、驢和營中一切的牲畜所遭的災殃與那災殃一樣。
ZECH|14|16|上來攻擊 耶路撒冷 的列國中所有剩下的人，要年年上來敬拜大君王－萬軍之耶和華，並守住棚節。
ZECH|14|17|地上萬族中，凡不上 耶路撒冷 敬拜大君王－萬軍之耶和華的，雨必不降在他們的地上。
ZECH|14|18|埃及 族若不上來，雨必不降在他們的地上；凡不上來守住棚節的列國，耶和華必用這災攻擊他們。
ZECH|14|19|這就是 埃及 的懲罰和那些不上來守住棚節之列國的懲罰。
ZECH|14|20|在那日，馬的鈴鐺上要刻上「歸耶和華為聖」。耶和華殿內的鍋必如祭壇前的碗一樣。
ZECH|14|21|耶路撒冷 和 猶大 一切的鍋都必歸萬軍之耶和華為聖。凡獻祭的都必來取這鍋，在其中煮肉。當那日，在萬軍之耶和華的殿中必不再有做買賣的人 。
