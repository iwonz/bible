ISA|1|1|The vision concerning Judah and Jerusalem that Isaiah son of Amoz saw during the reigns of Uzziah, Jotham, Ahaz and Hezekiah, kings of Judah.
ISA|1|2|Hear, O heavens! Listen, O earth! For the LORD has spoken: "I reared children and brought them up, but they have rebelled against me.
ISA|1|3|The ox knows his master, the donkey his owner's manger, but Israel does not know, my people do not understand."
ISA|1|4|Ah, sinful nation, a people loaded with guilt, a brood of evildoers, children given to corruption! They have forsaken the LORD; they have spurned the Holy One of Israel and turned their backs on him.
ISA|1|5|Why should you be beaten anymore? Why do you persist in rebellion? Your whole head is injured, your whole heart afflicted.
ISA|1|6|From the sole of your foot to the top of your head there is no soundness- only wounds and welts and open sores, not cleansed or bandaged or soothed with oil.
ISA|1|7|Your country is desolate, your cities burned with fire; your fields are being stripped by foreigners right before you, laid waste as when overthrown by strangers.
ISA|1|8|The Daughter of Zion is left like a shelter in a vineyard, like a hut in a field of melons, like a city under siege.
ISA|1|9|Unless the LORD Almighty had left us some survivors, we would have become like Sodom, we would have been like Gomorrah.
ISA|1|10|Hear the word of the LORD, you rulers of Sodom; listen to the law of our God, you people of Gomorrah!
ISA|1|11|"The multitude of your sacrifices- what are they to me?" says the LORD. "I have more than enough of burnt offerings, of rams and the fat of fattened animals; I have no pleasure in the blood of bulls and lambs and goats.
ISA|1|12|When you come to appear before me, who has asked this of you, this trampling of my courts?
ISA|1|13|Stop bringing meaningless offerings! Your incense is detestable to me. New Moons, Sabbaths and convocations- I cannot bear your evil assemblies.
ISA|1|14|Your New Moon festivals and your appointed feasts my soul hates. They have become a burden to me; I am weary of bearing them.
ISA|1|15|When you spread out your hands in prayer, I will hide my eyes from you; even if you offer many prayers, I will not listen. Your hands are full of blood;
ISA|1|16|wash and make yourselves clean. Take your evil deeds out of my sight! Stop doing wrong,
ISA|1|17|learn to do right! Seek justice, encourage the oppressed. Defend the cause of the fatherless, plead the case of the widow.
ISA|1|18|"Come now, let us reason together," says the LORD. "Though your sins are like scarlet, they shall be as white as snow; though they are red as crimson, they shall be like wool.
ISA|1|19|If you are willing and obedient, you will eat the best from the land;
ISA|1|20|but if you resist and rebel, you will be devoured by the sword." For the mouth of the LORD has spoken.
ISA|1|21|See how the faithful city has become a harlot! She once was full of justice; righteousness used to dwell in her- but now murderers!
ISA|1|22|Your silver has become dross, your choice wine is diluted with water.
ISA|1|23|Your rulers are rebels, companions of thieves; they all love bribes and chase after gifts. They do not defend the cause of the fatherless; the widow's case does not come before them.
ISA|1|24|Therefore the Lord, the LORD Almighty, the Mighty One of Israel, declares: "Ah, I will get relief from my foes and avenge myself on my enemies.
ISA|1|25|I will turn my hand against you; I will thoroughly purge away your dross and remove all your impurities.
ISA|1|26|I will restore your judges as in days of old, your counselors as at the beginning. Afterward you will be called the City of Righteousness, the Faithful City."
ISA|1|27|Zion will be redeemed with justice, her penitent ones with righteousness.
ISA|1|28|But rebels and sinners will both be broken, and those who forsake the LORD will perish.
ISA|1|29|"You will be ashamed because of the sacred oaks in which you have delighted; you will be disgraced because of the gardens that you have chosen.
ISA|1|30|You will be like an oak with fading leaves, like a garden without water.
ISA|1|31|The mighty man will become tinder and his work a spark; both will burn together, with no one to quench the fire."
ISA|2|1|This is what Isaiah son of Amoz saw concerning Judah and Jerusalem:
ISA|2|2|In the last days the mountain of the LORD's temple will be established as chief among the mountains; it will be raised above the hills, and all nations will stream to it.
ISA|2|3|Many peoples will come and say, "Come, let us go up to the mountain of the LORD, to the house of the God of Jacob. He will teach us his ways, so that we may walk in his paths." The law will go out from Zion, the word of the LORD from Jerusalem.
ISA|2|4|He will judge between the nations and will settle disputes for many peoples. They will beat their swords into plowshares and their spears into pruning hooks. Nation will not take up sword against nation, nor will they train for war anymore.
ISA|2|5|Come, O house of Jacob, let us walk in the light of the LORD.
ISA|2|6|You have abandoned your people, the house of Jacob. They are full of superstitions from the East; they practice divination like the Philistines and clasp hands with pagans.
ISA|2|7|Their land is full of silver and gold; there is no end to their treasures. Their land is full of horses; there is no end to their chariots.
ISA|2|8|Their land is full of idols; they bow down to the work of their hands, to what their fingers have made.
ISA|2|9|So man will be brought low and mankind humbled- do not forgive them.
ISA|2|10|Go into the rocks, hide in the ground from dread of the LORD and the splendor of his majesty!
ISA|2|11|The eyes of the arrogant man will be humbled and the pride of men brought low; the LORD alone will be exalted in that day.
ISA|2|12|The LORD Almighty has a day in store for all the proud and lofty, for all that is exalted (and they will be humbled),
ISA|2|13|for all the cedars of Lebanon, tall and lofty, and all the oaks of Bashan,
ISA|2|14|for all the towering mountains and all the high hills,
ISA|2|15|for every lofty tower and every fortified wall,
ISA|2|16|for every trading ship and every stately vessel.
ISA|2|17|The arrogance of man will be brought low and the pride of men humbled; the LORD alone will be exalted in that day,
ISA|2|18|and the idols will totally disappear.
ISA|2|19|Men will flee to caves in the rocks and to holes in the ground from dread of the LORD and the splendor of his majesty, when he rises to shake the earth.
ISA|2|20|In that day men will throw away to the rodents and bats their idols of silver and idols of gold, which they made to worship.
ISA|2|21|They will flee to caverns in the rocks and to the overhanging crags from dread of the LORD and the splendor of his majesty, when he rises to shake the earth.
ISA|2|22|Stop trusting in man, who has but a breath in his nostrils. Of what account is he?
ISA|3|1|See now, the Lord, the LORD Almighty, is about to take from Jerusalem and Judah both supply and support: all supplies of food and all supplies of water,
ISA|3|2|the hero and warrior, the judge and prophet, the soothsayer and elder,
ISA|3|3|the captain of fifty and man of rank, the counselor, skilled craftsman and clever enchanter.
ISA|3|4|I will make boys their officials; mere children will govern them.
ISA|3|5|People will oppress each other- man against man, neighbor against neighbor. The young will rise up against the old, the base against the honorable.
ISA|3|6|A man will seize one of his brothers at his father's home, and say, "You have a cloak, you be our leader; take charge of this heap of ruins!"
ISA|3|7|But in that day he will cry out, "I have no remedy. I have no food or clothing in my house; do not make me the leader of the people."
ISA|3|8|Jerusalem staggers, Judah is falling; their words and deeds are against the LORD, defying his glorious presence.
ISA|3|9|The look on their faces testifies against them; they parade their sin like Sodom; they do not hide it. Woe to them! They have brought disaster upon themselves.
ISA|3|10|Tell the righteous it will be well with them, for they will enjoy the fruit of their deeds.
ISA|3|11|Woe to the wicked! Disaster is upon them! They will be paid back for what their hands have done.
ISA|3|12|Youths oppress my people, women rule over them. O my people, your guides lead you astray; they turn you from the path.
ISA|3|13|The LORD takes his place in court; he rises to judge the people.
ISA|3|14|The LORD enters into judgment against the elders and leaders of his people: "It is you who have ruined my vineyard; the plunder from the poor is in your houses.
ISA|3|15|What do you mean by crushing my people and grinding the faces of the poor?" declares the Lord, the LORD Almighty.
ISA|3|16|The LORD says, "The women of Zion are haughty, walking along with outstretched necks, flirting with their eyes, tripping along with mincing steps, with ornaments jingling on their ankles.
ISA|3|17|Therefore the Lord will bring sores on the heads of the women of Zion; the LORD will make their scalps bald."
ISA|3|18|In that day the Lord will snatch away their finery: the bangles and headbands and crescent necklaces,
ISA|3|19|the earrings and bracelets and veils,
ISA|3|20|the headdresses and ankle chains and sashes, the perfume bottles and charms,
ISA|3|21|the signet rings and nose rings,
ISA|3|22|the fine robes and the capes and cloaks, the purses
ISA|3|23|and mirrors, and the linen garments and tiaras and shawls.
ISA|3|24|Instead of fragrance there will be a stench; instead of a sash, a rope; instead of well-dressed hair, baldness; instead of fine clothing, sackcloth; instead of beauty, branding.
ISA|3|25|Your men will fall by the sword, your warriors in battle.
ISA|3|26|The gates of Zion will lament and mourn; destitute, she will sit on the ground.
ISA|4|1|In that day seven women will take hold of one man and say, "We will eat our own food and provide our own clothes; only let us be called by your name. Take away our disgrace!"
ISA|4|2|In that day the Branch of the LORD will be beautiful and glorious, and the fruit of the land will be the pride and glory of the survivors in Israel.
ISA|4|3|Those who are left in Zion, who remain in Jerusalem, will be called holy, all who are recorded among the living in Jerusalem.
ISA|4|4|The Lord will wash away the filth of the women of Zion; he will cleanse the bloodstains from Jerusalem by a spirit of judgment and a spirit of fire.
ISA|4|5|Then the LORD will create over all of Mount Zion and over those who assemble there a cloud of smoke by day and a glow of flaming fire by night; over all the glory will be a canopy.
ISA|4|6|It will be a shelter and shade from the heat of the day, and a refuge and hiding place from the storm and rain.
ISA|5|1|I will sing for the one I love a song about his vineyard: My loved one had a vineyard on a fertile hillside.
ISA|5|2|He dug it up and cleared it of stones and planted it with the choicest vines. He built a watchtower in it and cut out a winepress as well. Then he looked for a crop of good grapes, but it yielded only bad fruit.
ISA|5|3|"Now you dwellers in Jerusalem and men of Judah, judge between me and my vineyard.
ISA|5|4|What more could have been done for my vineyard than I have done for it? When I looked for good grapes, why did it yield only bad?
ISA|5|5|Now I will tell you what I am going to do to my vineyard: I will take away its hedge, and it will be destroyed; I will break down its wall, and it will be trampled.
ISA|5|6|I will make it a wasteland, neither pruned nor cultivated, and briers and thorns will grow there. I will command the clouds not to rain on it."
ISA|5|7|The vineyard of the LORD Almighty is the house of Israel, and the men of Judah are the garden of his delight. And he looked for justice, but saw bloodshed; for righteousness, but heard cries of distress.
ISA|5|8|Woe to you who add house to house and join field to field till no space is left and you live alone in the land.
ISA|5|9|The LORD Almighty has declared in my hearing: "Surely the great houses will become desolate, the fine mansions left without occupants.
ISA|5|10|A ten-acre vineyard will produce only a bath of wine, a homer of seed only an ephah of grain."
ISA|5|11|Woe to those who rise early in the morning to run after their drinks, who stay up late at night till they are inflamed with wine.
ISA|5|12|They have harps and lyres at their banquets, tambourines and flutes and wine, but they have no regard for the deeds of the LORD, no respect for the work of his hands.
ISA|5|13|Therefore my people will go into exile for lack of understanding; their men of rank will die of hunger and their masses will be parched with thirst.
ISA|5|14|Therefore the grave enlarges its appetite and opens its mouth without limit; into it will descend their nobles and masses with all their brawlers and revelers.
ISA|5|15|So man will be brought low and mankind humbled, the eyes of the arrogant humbled.
ISA|5|16|But the LORD Almighty will be exalted by his justice, and the holy God will show himself holy by his righteousness.
ISA|5|17|Then sheep will graze as in their own pasture; lambs will feed among the ruins of the rich.
ISA|5|18|Woe to those who draw sin along with cords of deceit, and wickedness as with cart ropes,
ISA|5|19|to those who say, "Let God hurry, let him hasten his work so we may see it. Let it approach, let the plan of the Holy One of Israel come, so we may know it."
ISA|5|20|Woe to those who call evil good and good evil, who put darkness for light and light for darkness, who put bitter for sweet and sweet for bitter.
ISA|5|21|Woe to those who are wise in their own eyes and clever in their own sight.
ISA|5|22|Woe to those who are heroes at drinking wine and champions at mixing drinks,
ISA|5|23|who acquit the guilty for a bribe, but deny justice to the innocent.
ISA|5|24|Therefore, as tongues of fire lick up straw and as dry grass sinks down in the flames, so their roots will decay and their flowers blow away like dust; for they have rejected the law of the LORD Almighty and spurned the word of the Holy One of Israel.
ISA|5|25|Therefore the LORD's anger burns against his people; his hand is raised and he strikes them down. The mountains shake, and the dead bodies are like refuse in the streets. Yet for all this, his anger is not turned away, his hand is still upraised.
ISA|5|26|He lifts up a banner for the distant nations, he whistles for those at the ends of the earth. Here they come, swiftly and speedily!
ISA|5|27|Not one of them grows tired or stumbles, not one slumbers or sleeps; not a belt is loosened at the waist, not a sandal thong is broken.
ISA|5|28|Their arrows are sharp, all their bows are strung; their horses' hoofs seem like flint, their chariot wheels like a whirlwind.
ISA|5|29|Their roar is like that of the lion, they roar like young lions; they growl as they seize their prey and carry it off with no one to rescue.
ISA|5|30|In that day they will roar over it like the roaring of the sea. And if one looks at the land, he will see darkness and distress; even the light will be darkened by the clouds.
ISA|6|1|In the year that King Uzziah died, I saw the Lord seated on a throne, high and exalted, and the train of his robe filled the temple.
ISA|6|2|Above him were seraphs, each with six wings: With two wings they covered their faces, with two they covered their feet, and with two they were flying.
ISA|6|3|And they were calling to one another: "Holy, holy, holy is the LORD Almighty; the whole earth is full of his glory."
ISA|6|4|At the sound of their voices the doorposts and thresholds shook and the temple was filled with smoke.
ISA|6|5|"Woe to me!" I cried. "I am ruined! For I am a man of unclean lips, and I live among a people of unclean lips, and my eyes have seen the King, the LORD Almighty."
ISA|6|6|Then one of the seraphs flew to me with a live coal in his hand, which he had taken with tongs from the altar.
ISA|6|7|With it he touched my mouth and said, "See, this has touched your lips; your guilt is taken away and your sin atoned for."
ISA|6|8|Then I heard the voice of the Lord saying, "Whom shall I send? And who will go for us?" And I said, "Here am I. Send me!"
ISA|6|9|He said, "Go and tell this people: "'Be ever hearing, but never understanding; be ever seeing, but never perceiving.'
ISA|6|10|Make the heart of this people calloused; make their ears dull and close their eyes. Otherwise they might see with their eyes, hear with their ears, understand with their hearts, and turn and be healed."
ISA|6|11|Then I said, "For how long, O Lord?" And he answered: "Until the cities lie ruined and without inhabitant, until the houses are left deserted and the fields ruined and ravaged,
ISA|6|12|until the LORD has sent everyone far away and the land is utterly forsaken.
ISA|6|13|And though a tenth remains in the land, it will again be laid waste. But as the terebinth and oak leave stumps when they are cut down, so the holy seed will be the stump in the land."
ISA|7|1|When Ahaz son of Jotham, the son of Uzziah, was king of Judah, King Rezin of Aram and Pekah son of Remaliah king of Israel marched up to fight against Jerusalem, but they could not overpower it.
ISA|7|2|Now the house of David was told, "Aram has allied itself with Ephraim"; so the hearts of Ahaz and his people were shaken, as the trees of the forest are shaken by the wind.
ISA|7|3|Then the LORD said to Isaiah, "Go out, you and your son Shear-Jashub, to meet Ahaz at the end of the aqueduct of the Upper Pool, on the road to the Washerman's Field.
ISA|7|4|Say to him, 'Be careful, keep calm and don't be afraid. Do not lose heart because of these two smoldering stubs of firewood-because of the fierce anger of Rezin and Aram and of the son of Remaliah.
ISA|7|5|Aram, Ephraim and Remaliah's son have plotted your ruin, saying,
ISA|7|6|"Let us invade Judah; let us tear it apart and divide it among ourselves, and make the son of Tabeel king over it."
ISA|7|7|Yet this is what the Sovereign LORD says: "'It will not take place, it will not happen,
ISA|7|8|for the head of Aram is Damascus, and the head of Damascus is only Rezin. Within sixty-five years Ephraim will be too shattered to be a people.
ISA|7|9|The head of Ephraim is Samaria, and the head of Samaria is only Remaliah's son. If you do not stand firm in your faith, you will not stand at all.'"
ISA|7|10|Again the LORD spoke to Ahaz,
ISA|7|11|"Ask the LORD your God for a sign, whether in the deepest depths or in the highest heights."
ISA|7|12|But Ahaz said, "I will not ask; I will not put the LORD to the test."
ISA|7|13|Then Isaiah said, "Hear now, you house of David! Is it not enough to try the patience of men? Will you try the patience of my God also?
ISA|7|14|Therefore the Lord himself will give you a sign: The virgin will be with child and will give birth to a son, and will call him Immanuel.
ISA|7|15|He will eat curds and honey when he knows enough to reject the wrong and choose the right.
ISA|7|16|But before the boy knows enough to reject the wrong and choose the right, the land of the two kings you dread will be laid waste.
ISA|7|17|The LORD will bring on you and on your people and on the house of your father a time unlike any since Ephraim broke away from Judah-he will bring the king of Assyria."
ISA|7|18|In that day the LORD will whistle for flies from the distant streams of Egypt and for bees from the land of Assyria.
ISA|7|19|They will all come and settle in the steep ravines and in the crevices in the rocks, on all the thornbushes and at all the water holes.
ISA|7|20|In that day the Lord will use a razor hired from beyond the River -the king of Assyria-to shave your head and the hair of your legs, and to take off your beards also.
ISA|7|21|In that day, a man will keep alive a young cow and two goats.
ISA|7|22|And because of the abundance of the milk they give, he will have curds to eat. All who remain in the land will eat curds and honey.
ISA|7|23|In that day, in every place where there were a thousand vines worth a thousand silver shekels, there will be only briers and thorns.
ISA|7|24|Men will go there with bow and arrow, for the land will be covered with briers and thorns.
ISA|7|25|As for all the hills once cultivated by the hoe, you will no longer go there for fear of the briers and thorns; they will become places where cattle are turned loose and where sheep run.
ISA|8|1|The LORD said to me, "Take a large scroll and write on it with an ordinary pen: Maher-Shalal-Hash-Baz.
ISA|8|2|And I will call in Uriah the priest and Zechariah son of Jeberekiah as reliable witnesses for me."
ISA|8|3|Then I went to the prophetess, and she conceived and gave birth to a son. And the LORD said to me, "Name him Maher-Shalal-Hash-Baz.
ISA|8|4|Before the boy knows how to say 'My father' or 'My mother,' the wealth of Damascus and the plunder of Samaria will be carried off by the king of Assyria."
ISA|8|5|The LORD spoke to me again:
ISA|8|6|"Because this people has rejected the gently flowing waters of Shiloah and rejoices over Rezin and the son of Remaliah,
ISA|8|7|therefore the Lord is about to bring against them the mighty floodwaters of the River - the king of Assyria with all his pomp. It will overflow all its channels, run over all its banks
ISA|8|8|and sweep on into Judah, swirling over it, passing through it and reaching up to the neck. Its outspread wings will cover the breadth of your land, O Immanuel!"
ISA|8|9|Raise the war cry, you nations, and be shattered! Listen, all you distant lands. Prepare for battle, and be shattered! Prepare for battle, and be shattered!
ISA|8|10|Devise your strategy, but it will be thwarted; propose your plan, but it will not stand, for God is with us.
ISA|8|11|The LORD spoke to me with his strong hand upon me, warning me not to follow the way of this people. He said:
ISA|8|12|"Do not call conspiracy everything that these people call conspiracy; do not fear what they fear, and do not dread it.
ISA|8|13|The LORD Almighty is the one you are to regard as holy, he is the one you are to fear, he is the one you are to dread,
ISA|8|14|and he will be a sanctuary; but for both houses of Israel he will be a stone that causes men to stumble and a rock that makes them fall. And for the people of Jerusalem he will be a trap and a snare.
ISA|8|15|Many of them will stumble; they will fall and be broken, they will be snared and captured."
ISA|8|16|Bind up the testimony and seal up the law among my disciples.
ISA|8|17|I will wait for the LORD, who is hiding his face from the house of Jacob. I will put my trust in him.
ISA|8|18|Here am I, and the children the LORD has given me. We are signs and symbols in Israel from the LORD Almighty, who dwells on Mount Zion.
ISA|8|19|When men tell you to consult mediums and spiritists, who whisper and mutter, should not a people inquire of their God? Why consult the dead on behalf of the living?
ISA|8|20|To the law and to the testimony! If they do not speak according to this word, they have no light of dawn.
ISA|8|21|Distressed and hungry, they will roam through the land; when they are famished, they will become enraged and, looking upward, will curse their king and their God.
ISA|8|22|Then they will look toward the earth and see only distress and darkness and fearful gloom, and they will be thrust into utter darkness.
ISA|9|1|Nevertheless, there will be no more gloom for those who were in distress. In the past he humbled the land of Zebulun and the land of Naphtali, but in the future he will honor Galilee of the Gentiles, by the way of the sea, along the Jordan-
ISA|9|2|The people walking in darkness have seen a great light; on those living in the land of the shadow of death a light has dawned.
ISA|9|3|You have enlarged the nation and increased their joy; they rejoice before you as people rejoice at the harvest, as men rejoice when dividing the plunder.
ISA|9|4|For as in the day of Midian's defeat, you have shattered the yoke that burdens them, the bar across their shoulders, the rod of their oppressor.
ISA|9|5|Every warrior's boot used in battle and every garment rolled in blood will be destined for burning, will be fuel for the fire.
ISA|9|6|For to us a child is born, to us a son is given, and the government will be on his shoulders. And he will be called Wonderful Counselor, Mighty God, Everlasting Father, Prince of Peace.
ISA|9|7|Of the increase of his government and peace there will be no end. He will reign on David's throne and over his kingdom, establishing and upholding it with justice and righteousness from that time on and forever. The zeal of the LORD Almighty will accomplish this.
ISA|9|8|The Lord has sent a message against Jacob; it will fall on Israel.
ISA|9|9|All the people will know it- Ephraim and the inhabitants of Samaria- who say with pride and arrogance of heart,
ISA|9|10|"The bricks have fallen down, but we will rebuild with dressed stone; the fig trees have been felled, but we will replace them with cedars."
ISA|9|11|But the LORD has strengthened Rezin's foes against them and has spurred their enemies on.
ISA|9|12|Arameans from the east and Philistines from the west have devoured Israel with open mouth. Yet for all this, his anger is not turned away, his hand is still upraised.
ISA|9|13|But the people have not returned to him who struck them, nor have they sought the LORD Almighty.
ISA|9|14|So the LORD will cut off from Israel both head and tail, both palm branch and reed in a single day;
ISA|9|15|the elders and prominent men are the head, the prophets who teach lies are the tail.
ISA|9|16|Those who guide this people mislead them, and those who are guided are led astray.
ISA|9|17|Therefore the Lord will take no pleasure in the young men, nor will he pity the fatherless and widows, for everyone is ungodly and wicked, every mouth speaks vileness. Yet for all this, his anger is not turned away, his hand is still upraised.
ISA|9|18|Surely wickedness burns like a fire; it consumes briers and thorns, it sets the forest thickets ablaze, so that it rolls upward in a column of smoke.
ISA|9|19|By the wrath of the LORD Almighty the land will be scorched and the people will be fuel for the fire; no one will spare his brother.
ISA|9|20|On the right they will devour, but still be hungry; on the left they will eat, but not be satisfied. Each will feed on the flesh of his own offspring:
ISA|9|21|Manasseh will feed on Ephraim, and Ephraim on Manasseh; together they will turn against Judah. Yet for all this, his anger is not turned away, his hand is still upraised.
ISA|10|1|Woe to those who make unjust laws, to those who issue oppressive decrees,
ISA|10|2|to deprive the poor of their rights and withhold justice from the oppressed of my people, making widows their prey and robbing the fatherless.
ISA|10|3|What will you do on the day of reckoning, when disaster comes from afar? To whom will you run for help? Where will you leave your riches?
ISA|10|4|Nothing will remain but to cringe among the captives or fall among the slain. Yet for all this, his anger is not turned away, his hand is still upraised.
ISA|10|5|"Woe to the Assyrian, the rod of my anger, in whose hand is the club of my wrath!
ISA|10|6|I send him against a godless nation, I dispatch him against a people who anger me, to seize loot and snatch plunder, and to trample them down like mud in the streets.
ISA|10|7|But this is not what he intends, this is not what he has in mind; his purpose is to destroy, to put an end to many nations.
ISA|10|8|'Are not my commanders all kings?' he says.
ISA|10|9|'Has not Calno fared like Carchemish? Is not Hamath like Arpad, and Samaria like Damascus?
ISA|10|10|As my hand seized the kingdoms of the idols, kingdoms whose images excelled those of Jerusalem and Samaria-
ISA|10|11|shall I not deal with Jerusalem and her images as I dealt with Samaria and her idols?'"
ISA|10|12|When the Lord has finished all his work against Mount Zion and Jerusalem, he will say, "I will punish the king of Assyria for the willful pride of his heart and the haughty look in his eyes.
ISA|10|13|For he says: "'By the strength of my hand I have done this, and by my wisdom, because I have understanding. I removed the boundaries of nations, I plundered their treasures; like a mighty one I subdued their kings.
ISA|10|14|As one reaches into a nest, so my hand reached for the wealth of the nations; as men gather abandoned eggs, so I gathered all the countries; not one flapped a wing, or opened its mouth to chirp.'"
ISA|10|15|Does the ax raise itself above him who swings it, or the saw boast against him who uses it? As if a rod were to wield him who lifts it up, or a club brandish him who is not wood!
ISA|10|16|Therefore, the Lord, the LORD Almighty, will send a wasting disease upon his sturdy warriors; under his pomp a fire will be kindled like a blazing flame.
ISA|10|17|The Light of Israel will become a fire, their Holy One a flame; in a single day it will burn and consume his thorns and his briers.
ISA|10|18|The splendor of his forests and fertile fields it will completely destroy, as when a sick man wastes away.
ISA|10|19|And the remaining trees of his forests will be so few that a child could write them down.
ISA|10|20|In that day the remnant of Israel, the survivors of the house of Jacob, will no longer rely on him who struck them down but will truly rely on the LORD, the Holy One of Israel.
ISA|10|21|A remnant will return, a remnant of Jacob will return to the Mighty God.
ISA|10|22|Though your people, O Israel, be like the sand by the sea, only a remnant will return. Destruction has been decreed, overwhelming and righteous.
ISA|10|23|The Lord, the LORD Almighty, will carry out the destruction decreed upon the whole land.
ISA|10|24|Therefore, this is what the Lord, the LORD Almighty, says: "O my people who live in Zion, do not be afraid of the Assyrians, who beat you with a rod and lift up a club against you, as Egypt did.
ISA|10|25|Very soon my anger against you will end and my wrath will be directed to their destruction."
ISA|10|26|The LORD Almighty will lash them with a whip, as when he struck down Midian at the rock of Oreb; and he will raise his staff over the waters, as he did in Egypt.
ISA|10|27|In that day their burden will be lifted from your shoulders, their yoke from your neck; the yoke will be broken because you have grown so fat.
ISA|10|28|They enter Aiath; they pass through Migron; they store supplies at Micmash.
ISA|10|29|They go over the pass, and say, "We will camp overnight at Geba." Ramah trembles; Gibeah of Saul flees.
ISA|10|30|Cry out, O Daughter of Gallim! Listen, O Laishah! Poor Anathoth!
ISA|10|31|Madmenah is in flight; the people of Gebim take cover.
ISA|10|32|This day they will halt at Nob; they will shake their fist at the mount of the Daughter of Zion, at the hill of Jerusalem.
ISA|10|33|See, the Lord, the LORD Almighty, will lop off the boughs with great power. The lofty trees will be felled, the tall ones will be brought low.
ISA|10|34|He will cut down the forest thickets with an ax; Lebanon will fall before the Mighty One.
ISA|11|1|A shoot will come up from the stump of Jesse; from his roots a Branch will bear fruit.
ISA|11|2|The Spirit of the LORD will rest on him- the Spirit of wisdom and of understanding, the Spirit of counsel and of power, the Spirit of knowledge and of the fear of the LORD -
ISA|11|3|and he will delight in the fear of the LORD. He will not judge by what he sees with his eyes, or decide by what he hears with his ears;
ISA|11|4|but with righteousness he will judge the needy, with justice he will give decisions for the poor of the earth. He will strike the earth with the rod of his mouth; with the breath of his lips he will slay the wicked.
ISA|11|5|Righteousness will be his belt and faithfulness the sash around his waist.
ISA|11|6|The wolf will live with the lamb, the leopard will lie down with the goat, the calf and the lion and the yearling together; and a little child will lead them.
ISA|11|7|The cow will feed with the bear, their young will lie down together, and the lion will eat straw like the ox.
ISA|11|8|The infant will play near the hole of the cobra, and the young child put his hand into the viper's nest.
ISA|11|9|They will neither harm nor destroy on all my holy mountain, for the earth will be full of the knowledge of the LORD as the waters cover the sea.
ISA|11|10|In that day the Root of Jesse will stand as a banner for the peoples; the nations will rally to him, and his place of rest will be glorious.
ISA|11|11|In that day the Lord will reach out his hand a second time to reclaim the remnant that is left of his people from Assyria, from Lower Egypt, from Upper Egypt, from Cush, from Elam, from Babylonia, from Hamath and from the islands of the sea.
ISA|11|12|He will raise a banner for the nations and gather the exiles of Israel; he will assemble the scattered people of Judah from the four quarters of the earth.
ISA|11|13|Ephraim's jealousy will vanish, and Judah's enemies will be cut off; Ephraim will not be jealous of Judah, nor Judah hostile toward Ephraim.
ISA|11|14|They will swoop down on the slopes of Philistia to the west; together they will plunder the people to the east. They will lay hands on Edom and Moab, and the Ammonites will be subject to them.
ISA|11|15|The LORD will dry up the gulf of the Egyptian sea; with a scorching wind he will sweep his hand over the Euphrates River. He will break it up into seven streams so that men can cross over in sandals.
ISA|11|16|There will be a highway for the remnant of his people that is left from Assyria, as there was for Israel when they came up from Egypt.
ISA|12|1|In that day you will say: "I will praise you, O LORD. Although you were angry with me, your anger has turned away and you have comforted me.
ISA|12|2|Surely God is my salvation; I will trust and not be afraid. The LORD, the LORD, is my strength and my song; he has become my salvation."
ISA|12|3|With joy you will draw water from the wells of salvation.
ISA|12|4|In that day you will say: "Give thanks to the LORD, call on his name; make known among the nations what he has done, and proclaim that his name is exalted.
ISA|12|5|Sing to the LORD, for he has done glorious things; let this be known to all the world.
ISA|12|6|Shout aloud and sing for joy, people of Zion, for great is the Holy One of Israel among you."
ISA|13|1|An oracle concerning Babylon that Isaiah son of Amoz saw:
ISA|13|2|Raise a banner on a bare hilltop, shout to them; beckon to them to enter the gates of the nobles.
ISA|13|3|I have commanded my holy ones; I have summoned my warriors to carry out my wrath- those who rejoice in my triumph.
ISA|13|4|Listen, a noise on the mountains, like that of a great multitude! Listen, an uproar among the kingdoms, like nations massing together! The LORD Almighty is mustering an army for war.
ISA|13|5|They come from faraway lands, from the ends of the heavens- the LORD and the weapons of his wrath- to destroy the whole country.
ISA|13|6|Wail, for the day of the LORD is near; it will come like destruction from the Almighty.
ISA|13|7|Because of this, all hands will go limp, every man's heart will melt.
ISA|13|8|Terror will seize them, pain and anguish will grip them; they will writhe like a woman in labor. They will look aghast at each other, their faces aflame.
ISA|13|9|See, the day of the LORD is coming -a cruel day, with wrath and fierce anger- to make the land desolate and destroy the sinners within it.
ISA|13|10|The stars of heaven and their constellations will not show their light. The rising sun will be darkened and the moon will not give its light.
ISA|13|11|I will punish the world for its evil, the wicked for their sins. I will put an end to the arrogance of the haughty and will humble the pride of the ruthless.
ISA|13|12|I will make man scarcer than pure gold, more rare than the gold of Ophir.
ISA|13|13|Therefore I will make the heavens tremble; and the earth will shake from its place at the wrath of the LORD Almighty, in the day of his burning anger.
ISA|13|14|Like a hunted gazelle, like sheep without a shepherd, each will return to his own people, each will flee to his native land.
ISA|13|15|Whoever is captured will be thrust through; all who are caught will fall by the sword.
ISA|13|16|Their infants will be dashed to pieces before their eyes; their houses will be looted and their wives ravished.
ISA|13|17|See, I will stir up against them the Medes, who do not care for silver and have no delight in gold.
ISA|13|18|Their bows will strike down the young men; they will have no mercy on infants nor will they look with compassion on children.
ISA|13|19|Babylon, the jewel of kingdoms, the glory of the Babylonians' pride, will be overthrown by God like Sodom and Gomorrah.
ISA|13|20|She will never be inhabited or lived in through all generations; no Arab will pitch his tent there, no shepherd will rest his flocks there.
ISA|13|21|But desert creatures will lie there, jackals will fill her houses; there the owls will dwell, and there the wild goats will leap about.
ISA|13|22|Hyenas will howl in her strongholds, jackals in her luxurious palaces. Her time is at hand, and her days will not be prolonged.
ISA|14|1|The LORD will have compassion on Jacob; once again he will choose Israel and will settle them in their own land. Aliens will join them and unite with the house of Jacob.
ISA|14|2|Nations will take them and bring them to their own place. And the house of Israel will possess the nations as menservants and maidservants in the LORD's land. They will make captives of their captors and rule over their oppressors.
ISA|14|3|On the day the LORD gives you relief from suffering and turmoil and cruel bondage,
ISA|14|4|you will take up this taunt against the king of Babylon: How the oppressor has come to an end! How his fury has ended!
ISA|14|5|The LORD has broken the rod of the wicked, the scepter of the rulers,
ISA|14|6|which in anger struck down peoples with unceasing blows, and in fury subdued nations with relentless aggression.
ISA|14|7|All the lands are at rest and at peace; they break into singing.
ISA|14|8|Even the pine trees and the cedars of Lebanon exult over you and say, "Now that you have been laid low, no woodsman comes to cut us down."
ISA|14|9|The grave below is all astir to meet you at your coming; it rouses the spirits of the departed to greet you- all those who were leaders in the world; it makes them rise from their thrones- all those who were kings over the nations.
ISA|14|10|They will all respond, they will say to you, "You also have become weak, as we are; you have become like us."
ISA|14|11|All your pomp has been brought down to the grave, along with the noise of your harps; maggots are spread out beneath you and worms cover you.
ISA|14|12|How you have fallen from heaven, O morning star, son of the dawn! You have been cast down to the earth, you who once laid low the nations!
ISA|14|13|You said in your heart, "I will ascend to heaven; I will raise my throne above the stars of God; I will sit enthroned on the mount of assembly, on the utmost heights of the sacred mountain.
ISA|14|14|I will ascend above the tops of the clouds; I will make myself like the Most High."
ISA|14|15|But you are brought down to the grave, to the depths of the pit.
ISA|14|16|Those who see you stare at you, they ponder your fate: "Is this the man who shook the earth and made kingdoms tremble,
ISA|14|17|the man who made the world a desert, who overthrew its cities and would not let his captives go home?"
ISA|14|18|All the kings of the nations lie in state, each in his own tomb.
ISA|14|19|But you are cast out of your tomb like a rejected branch; you are covered with the slain, with those pierced by the sword, those who descend to the stones of the pit. Like a corpse trampled underfoot,
ISA|14|20|you will not join them in burial, for you have destroyed your land and killed your people. The offspring of the wicked will never be mentioned again.
ISA|14|21|Prepare a place to slaughter his sons for the sins of their forefathers; they are not to rise to inherit the land and cover the earth with their cities.
ISA|14|22|"I will rise up against them," declares the LORD Almighty. "I will cut off from Babylon her name and survivors, her offspring and descendants," declares the LORD.
ISA|14|23|"I will turn her into a place for owls and into swampland; I will sweep her with the broom of destruction," declares the LORD Almighty.
ISA|14|24|The LORD Almighty has sworn, "Surely, as I have planned, so it will be, and as I have purposed, so it will stand.
ISA|14|25|I will crush the Assyrian in my land; on my mountains I will trample him down. His yoke will be taken from my people, and his burden removed from their shoulders."
ISA|14|26|This is the plan determined for the whole world; this is the hand stretched out over all nations.
ISA|14|27|For the LORD Almighty has purposed, and who can thwart him? His hand is stretched out, and who can turn it back?
ISA|14|28|This oracle came in the year King Ahaz died:
ISA|14|29|Do not rejoice, all you Philistines, that the rod that struck you is broken; from the root of that snake will spring up a viper, its fruit will be a darting, venomous serpent.
ISA|14|30|The poorest of the poor will find pasture, and the needy will lie down in safety. But your root I will destroy by famine; it will slay your survivors.
ISA|14|31|Wail, O gate! Howl, O city! Melt away, all you Philistines! A cloud of smoke comes from the north, and there is not a straggler in its ranks.
ISA|14|32|What answer shall be given to the envoys of that nation? "The LORD has established Zion, and in her his afflicted people will find refuge."
ISA|15|1|An oracle concerning Moab: Ar in Moab is ruined, destroyed in a night! Kir in Moab is ruined, destroyed in a night!
ISA|15|2|Dibon goes up to its temple, to its high places to weep; Moab wails over Nebo and Medeba. Every head is shaved and every beard cut off.
ISA|15|3|In the streets they wear sackcloth; on the roofs and in the public squares they all wail, prostrate with weeping.
ISA|15|4|Heshbon and Elealeh cry out, their voices are heard all the way to Jahaz. Therefore the armed men of Moab cry out, and their hearts are faint.
ISA|15|5|My heart cries out over Moab; her fugitives flee as far as Zoar, as far as Eglath Shelishiyah. They go up the way to Luhith, weeping as they go; on the road to Horonaim they lament their destruction.
ISA|15|6|The waters of Nimrim are dried up and the grass is withered; the vegetation is gone and nothing green is left.
ISA|15|7|So the wealth they have acquired and stored up they carry away over the Ravine of the Poplars.
ISA|15|8|Their outcry echoes along the border of Moab; their wailing reaches as far as Eglaim, their lamentation as far as Beer Elim.
ISA|15|9|Dimon's waters are full of blood, but I will bring still more upon Dimon - a lion upon the fugitives of Moab and upon those who remain in the land.
ISA|16|1|Send lambs as tribute to the ruler of the land, from Sela, across the desert, to the mount of the Daughter of Zion.
ISA|16|2|Like fluttering birds pushed from the nest, so are the women of Moab at the fords of the Arnon.
ISA|16|3|"Give us counsel, render a decision. Make your shadow like night- at high noon. Hide the fugitives, do not betray the refugees.
ISA|16|4|Let the Moabite fugitives stay with you; be their shelter from the destroyer." The oppressor will come to an end, and destruction will cease; the aggressor will vanish from the land.
ISA|16|5|In love a throne will be established; in faithfulness a man will sit on it- one from the house of David- one who in judging seeks justice and speeds the cause of righteousness.
ISA|16|6|We have heard of Moab's pride- her overweening pride and conceit, her pride and her insolence- but her boasts are empty.
ISA|16|7|Therefore the Moabites wail, they wail together for Moab. Lament and grieve for the men of Kir Hareseth.
ISA|16|8|The fields of Heshbon wither, the vines of Sibmah also. The rulers of the nations have trampled down the choicest vines, which once reached Jazer and spread toward the desert. Their shoots spread out and went as far as the sea.
ISA|16|9|So I weep, as Jazer weeps, for the vines of Sibmah. O Heshbon, O Elealeh, I drench you with tears! The shouts of joy over your ripened fruit and over your harvests have been stilled.
ISA|16|10|Joy and gladness are taken away from the orchards; no one sings or shouts in the vineyards; no one treads out wine at the presses, for I have put an end to the shouting.
ISA|16|11|My heart laments for Moab like a harp, my inmost being for Kir Hareseth.
ISA|16|12|When Moab appears at her high place, she only wears herself out; when she goes to her shrine to pray, it is to no avail.
ISA|16|13|This is the word the LORD has already spoken concerning Moab.
ISA|16|14|But now the LORD says: "Within three years, as a servant bound by contract would count them, Moab's splendor and all her many people will be despised, and her survivors will be very few and feeble."
ISA|17|1|An oracle concerning Damascus: "See, Damascus will no longer be a city but will become a heap of ruins.
ISA|17|2|The cities of Aroer will be deserted and left to flocks, which will lie down, with no one to make them afraid.
ISA|17|3|The fortified city will disappear from Ephraim, and royal power from Damascus; the remnant of Aram will be like the glory of the Israelites," declares the LORD Almighty.
ISA|17|4|"In that day the glory of Jacob will fade; the fat of his body will waste away.
ISA|17|5|It will be as when a reaper gathers the standing grain and harvests the grain with his arm- as when a man gleans heads of grain in the Valley of Rephaim.
ISA|17|6|Yet some gleanings will remain, as when an olive tree is beaten, leaving two or three olives on the topmost branches, four or five on the fruitful boughs," declares the LORD, the God of Israel.
ISA|17|7|In that day men will look to their Maker and turn their eyes to the Holy One of Israel.
ISA|17|8|They will not look to the altars, the work of their hands, and they will have no regard for the Asherah poles and the incense altars their fingers have made.
ISA|17|9|In that day their strong cities, which they left because of the Israelites, will be like places abandoned to thickets and undergrowth. And all will be desolation.
ISA|17|10|You have forgotten God your Savior; you have not remembered the Rock, your fortress. Therefore, though you set out the finest plants and plant imported vines,
ISA|17|11|though on the day you set them out, you make them grow, and on the morning when you plant them, you bring them to bud, yet the harvest will be as nothing in the day of disease and incurable pain.
ISA|17|12|Oh, the raging of many nations- they rage like the raging sea! Oh, the uproar of the peoples- they roar like the roaring of great waters!
ISA|17|13|Although the peoples roar like the roar of surging waters, when he rebukes them they flee far away, driven before the wind like chaff on the hills, like tumbleweed before a gale.
ISA|17|14|In the evening, sudden terror! Before the morning, they are gone! This is the portion of those who loot us, the lot of those who plunder us.
ISA|18|1|Woe to the land of whirring wings along the rivers of Cush,
ISA|18|2|which sends envoys by sea in papyrus boats over the water. Go, swift messengers, to a people tall and smooth-skinned, to a people feared far and wide, an aggressive nation of strange speech, whose land is divided by rivers.
ISA|18|3|All you people of the world, you who live on the earth, when a banner is raised on the mountains, you will see it, and when a trumpet sounds, you will hear it.
ISA|18|4|This is what the LORD says to me: "I will remain quiet and will look on from my dwelling place, like shimmering heat in the sunshine, like a cloud of dew in the heat of harvest."
ISA|18|5|For, before the harvest, when the blossom is gone and the flower becomes a ripening grape, he will cut off the shoots with pruning knives, and cut down and take away the spreading branches.
ISA|18|6|They will all be left to the mountain birds of prey and to the wild animals; the birds will feed on them all summer, the wild animals all winter.
ISA|18|7|At that time gifts will be brought to the LORD Almighty from a people tall and smooth-skinned, from a people feared far and wide, an aggressive nation of strange speech, whose land is divided by rivers- the gifts will be brought to Mount Zion, the place of the Name of the LORD Almighty.
ISA|19|1|An oracle concerning Egypt: See, the LORD rides on a swift cloud and is coming to Egypt. The idols of Egypt tremble before him, and the hearts of the Egyptians melt within them.
ISA|19|2|"I will stir up Egyptian against Egyptian- brother will fight against brother, neighbor against neighbor, city against city, kingdom against kingdom.
ISA|19|3|The Egyptians will lose heart, and I will bring their plans to nothing; they will consult the idols and the spirits of the dead, the mediums and the spiritists.
ISA|19|4|I will hand the Egyptians over to the power of a cruel master, and a fierce king will rule over them," declares the Lord, the LORD Almighty.
ISA|19|5|The waters of the river will dry up, and the riverbed will be parched and dry.
ISA|19|6|The canals will stink; the streams of Egypt will dwindle and dry up. The reeds and rushes will wither,
ISA|19|7|also the plants along the Nile, at the mouth of the river. Every sown field along the Nile will become parched, will blow away and be no more.
ISA|19|8|The fishermen will groan and lament, all who cast hooks into the Nile; those who throw nets on the water will pine away.
ISA|19|9|Those who work with combed flax will despair, the weavers of fine linen will lose hope.
ISA|19|10|The workers in cloth will be dejected, and all the wage earners will be sick at heart.
ISA|19|11|The officials of Zoan are nothing but fools; the wise counselors of Pharaoh give senseless advice. How can you say to Pharaoh, "I am one of the wise men, a disciple of the ancient kings"?
ISA|19|12|Where are your wise men now? Let them show you and make known what the LORD Almighty has planned against Egypt.
ISA|19|13|The officials of Zoan have become fools, the leaders of Memphis are deceived; the cornerstones of her peoples have led Egypt astray.
ISA|19|14|The LORD has poured into them a spirit of dizziness; they make Egypt stagger in all that she does, as a drunkard staggers around in his vomit.
ISA|19|15|There is nothing Egypt can do- head or tail, palm branch or reed.
ISA|19|16|In that day the Egyptians will be like women. They will shudder with fear at the uplifted hand that the LORD Almighty raises against them.
ISA|19|17|And the land of Judah will bring terror to the Egyptians; everyone to whom Judah is mentioned will be terrified, because of what the LORD Almighty is planning against them.
ISA|19|18|In that day five cities in Egypt will speak the language of Canaan and swear allegiance to the LORD Almighty. One of them will be called the City of Destruction.
ISA|19|19|In that day there will be an altar to the LORD in the heart of Egypt, and a monument to the LORD at its border.
ISA|19|20|It will be a sign and witness to the LORD Almighty in the land of Egypt. When they cry out to the LORD because of their oppressors, he will send them a savior and defender, and he will rescue them.
ISA|19|21|So the LORD will make himself known to the Egyptians, and in that day they will acknowledge the LORD. They will worship with sacrifices and grain offerings; they will make vows to the LORD and keep them.
ISA|19|22|The LORD will strike Egypt with a plague; he will strike them and heal them. They will turn to the LORD, and he will respond to their pleas and heal them.
ISA|19|23|In that day there will be a highway from Egypt to Assyria. The Assyrians will go to Egypt and the Egyptians to Assyria. The Egyptians and Assyrians will worship together.
ISA|19|24|In that day Israel will be the third, along with Egypt and Assyria, a blessing on the earth.
ISA|19|25|The LORD Almighty will bless them, saying, "Blessed be Egypt my people, Assyria my handiwork, and Israel my inheritance."
ISA|20|1|In the year that the supreme commander, sent by Sargon king of Assyria, came to Ashdod and attacked and captured it-
ISA|20|2|at that time the LORD spoke through Isaiah son of Amoz. He said to him, "Take off the sackcloth from your body and the sandals from your feet." And he did so, going around stripped and barefoot.
ISA|20|3|Then the LORD said, "Just as my servant Isaiah has gone stripped and barefoot for three years, as a sign and portent against Egypt and Cush,
ISA|20|4|so the king of Assyria will lead away stripped and barefoot the Egyptian captives and Cushite exiles, young and old, with buttocks bared-to Egypt's shame.
ISA|20|5|Those who trusted in Cush and boasted in Egypt will be afraid and put to shame.
ISA|20|6|In that day the people who live on this coast will say, 'See what has happened to those we relied on, those we fled to for help and deliverance from the king of Assyria! How then can we escape?'"
ISA|21|1|An oracle concerning the Desert by the Sea: Like whirlwinds sweeping through the southland, an invader comes from the desert, from a land of terror.
ISA|21|2|A dire vision has been shown to me: The traitor betrays, the looter takes loot. Elam, attack! Media, lay siege! I will bring to an end all the groaning she caused.
ISA|21|3|At this my body is racked with pain, pangs seize me, like those of a woman in labor; I am staggered by what I hear, I am bewildered by what I see.
ISA|21|4|My heart falters, fear makes me tremble; the twilight I longed for has become a horror to me.
ISA|21|5|They set the tables, they spread the rugs, they eat, they drink! Get up, you officers, oil the shields!
ISA|21|6|This is what the Lord says to me: "Go, post a lookout and have him report what he sees.
ISA|21|7|When he sees chariots with teams of horses, riders on donkeys or riders on camels, let him be alert, fully alert."
ISA|21|8|And the lookout shouted, "Day after day, my lord, I stand on the watchtower; every night I stay at my post.
ISA|21|9|Look, here comes a man in a chariot with a team of horses. And he gives back the answer: 'Babylon has fallen, has fallen! All the images of its gods lie shattered on the ground!'"
ISA|21|10|O my people, crushed on the threshing floor, I tell you what I have heard from the LORD Almighty, from the God of Israel.
ISA|21|11|An oracle concerning Dumah: Someone calls to me from Seir, "Watchman, what is left of the night? Watchman, what is left of the night?"
ISA|21|12|The watchman replies, "Morning is coming, but also the night. If you would ask, then ask; and come back yet again."
ISA|21|13|An oracle concerning Arabia: You caravans of Dedanites, who camp in the thickets of Arabia,
ISA|21|14|bring water for the thirsty; you who live in Tema, bring food for the fugitives.
ISA|21|15|They flee from the sword, from the drawn sword, from the bent bow and from the heat of battle.
ISA|21|16|This is what the Lord says to me: "Within one year, as a servant bound by contract would count it, all the pomp of Kedar will come to an end.
ISA|21|17|The survivors of the bowmen, the warriors of Kedar, will be few." The LORD, the God of Israel, has spoken.
ISA|22|1|An oracle concerning the Valley of Vision: What troubles you now, that you have all gone up on the roofs,
ISA|22|2|O town full of commotion, O city of tumult and revelry? Your slain were not killed by the sword, nor did they die in battle.
ISA|22|3|All your leaders have fled together; they have been captured without using the bow. All you who were caught were taken prisoner together, having fled while the enemy was still far away.
ISA|22|4|Therefore I said, "Turn away from me; let me weep bitterly. Do not try to console me over the destruction of my people."
ISA|22|5|The Lord, the LORD Almighty, has a day of tumult and trampling and terror in the Valley of Vision, a day of battering down walls and of crying out to the mountains.
ISA|22|6|Elam takes up the quiver, with her charioteers and horses; Kir uncovers the shield.
ISA|22|7|Your choicest valleys are full of chariots, and horsemen are posted at the city gates;
ISA|22|8|the defenses of Judah are stripped away. And you looked in that day to the weapons in the Palace of the Forest;
ISA|22|9|you saw that the City of David had many breaches in its defenses; you stored up water in the Lower Pool.
ISA|22|10|You counted the buildings in Jerusalem and tore down houses to strengthen the wall.
ISA|22|11|You built a reservoir between the two walls for the water of the Old Pool, but you did not look to the One who made it, or have regard for the One who planned it long ago.
ISA|22|12|The Lord, the LORD Almighty, called you on that day to weep and to wail, to tear out your hair and put on sackcloth.
ISA|22|13|But see, there is joy and revelry, slaughtering of cattle and killing of sheep, eating of meat and drinking of wine! "Let us eat and drink," you say, "for tomorrow we die!"
ISA|22|14|The LORD Almighty has revealed this in my hearing: "Till your dying day this sin will not be atoned for," says the Lord, the LORD Almighty.
ISA|22|15|This is what the Lord, the LORD Almighty, says: "Go, say to this steward, to Shebna, who is in charge of the palace:
ISA|22|16|What are you doing here and who gave you permission to cut out a grave for yourself here, hewing your grave on the height and chiseling your resting place in the rock?
ISA|22|17|"Beware, the LORD is about to take firm hold of you and hurl you away, O you mighty man.
ISA|22|18|He will roll you up tightly like a ball and throw you into a large country. There you will die and there your splendid chariots will remain- you disgrace to your master's house!
ISA|22|19|I will depose you from your office, and you will be ousted from your position.
ISA|22|20|"In that day I will summon my servant, Eliakim son of Hilkiah.
ISA|22|21|I will clothe him with your robe and fasten your sash around him and hand your authority over to him. He will be a father to those who live in Jerusalem and to the house of Judah.
ISA|22|22|I will place on his shoulder the key to the house of David; what he opens no one can shut, and what he shuts no one can open.
ISA|22|23|I will drive him like a peg into a firm place; he will be a seat of honor for the house of his father.
ISA|22|24|All the glory of his family will hang on him: its offspring and offshoots-all its lesser vessels, from the bowls to all the jars.
ISA|22|25|"In that day," declares the LORD Almighty, "the peg driven into the firm place will give way; it will be sheared off and will fall, and the load hanging on it will be cut down." The LORD has spoken.
ISA|23|1|An oracle concerning Tyre: Wail, O ships of Tarshish! For Tyre is destroyed and left without house or harbor. From the land of Cyprus word has come to them.
ISA|23|2|Be silent, you people of the island and you merchants of Sidon, whom the seafarers have enriched.
ISA|23|3|On the great waters came the grain of the Shihor; the harvest of the Nile was the revenue of Tyre, and she became the marketplace of the nations.
ISA|23|4|Be ashamed, O Sidon, and you, O fortress of the sea, for the sea has spoken: "I have neither been in labor nor given birth; I have neither reared sons nor brought up daughters."
ISA|23|5|When word comes to Egypt, they will be in anguish at the report from Tyre.
ISA|23|6|Cross over to Tarshish; wail, you people of the island.
ISA|23|7|Is this your city of revelry, the old, old city, whose feet have taken her to settle in far-off lands?
ISA|23|8|Who planned this against Tyre, the bestower of crowns, whose merchants are princes, whose traders are renowned in the earth?
ISA|23|9|The LORD Almighty planned it, to bring low the pride of all glory and to humble all who are renowned on the earth.
ISA|23|10|Till your land as along the Nile, O Daughter of Tarshish, for you no longer have a harbor.
ISA|23|11|The LORD has stretched out his hand over the sea and made its kingdoms tremble. He has given an order concerning Phoenicia that her fortresses be destroyed.
ISA|23|12|He said, "No more of your reveling, O Virgin Daughter of Sidon, now crushed! "Up, cross over to Cyprus; even there you will find no rest."
ISA|23|13|Look at the land of the Babylonians, this people that is now of no account! The Assyrians have made it a place for desert creatures; they raised up their siege towers, they stripped its fortresses bare and turned it into a ruin.
ISA|23|14|Wail, you ships of Tarshish; your fortress is destroyed!
ISA|23|15|At that time Tyre will be forgotten for seventy years, the span of a king's life. But at the end of these seventy years, it will happen to Tyre as in the song of the prostitute:
ISA|23|16|"Take up a harp, walk through the city, O prostitute forgotten; play the harp well, sing many a song, so that you will be remembered."
ISA|23|17|At the end of seventy years, the LORD will deal with Tyre. She will return to her hire as a prostitute and will ply her trade with all the kingdoms on the face of the earth.
ISA|23|18|Yet her profit and her earnings will be set apart for the LORD; they will not be stored up or hoarded. Her profits will go to those who live before the LORD, for abundant food and fine clothes.
ISA|24|1|See, the LORD is going to lay waste the earth and devastate it; he will ruin its face and scatter its inhabitants-
ISA|24|2|it will be the same for priest as for people, for master as for servant, for mistress as for maid, for seller as for buyer, for borrower as for lender, for debtor as for creditor.
ISA|24|3|The earth will be completely laid waste and totally plundered. The LORD has spoken this word.
ISA|24|4|The earth dries up and withers, the world languishes and withers, the exalted of the earth languish.
ISA|24|5|The earth is defiled by its people; they have disobeyed the laws, violated the statutes and broken the everlasting covenant.
ISA|24|6|Therefore a curse consumes the earth; its people must bear their guilt. Therefore earth's inhabitants are burned up, and very few are left.
ISA|24|7|The new wine dries up and the vine withers; all the merrymakers groan.
ISA|24|8|The gaiety of the tambourines is stilled, the noise of the revelers has stopped, the joyful harp is silent.
ISA|24|9|No longer do they drink wine with a song; the beer is bitter to its drinkers.
ISA|24|10|The ruined city lies desolate; the entrance to every house is barred.
ISA|24|11|In the streets they cry out for wine; all joy turns to gloom, all gaiety is banished from the earth.
ISA|24|12|The city is left in ruins, its gate is battered to pieces.
ISA|24|13|So will it be on the earth and among the nations, as when an olive tree is beaten, or as when gleanings are left after the grape harvest.
ISA|24|14|They raise their voices, they shout for joy; from the west they acclaim the LORD's majesty.
ISA|24|15|Therefore in the east give glory to the LORD; exalt the name of the LORD, the God of Israel, in the islands of the sea.
ISA|24|16|From the ends of the earth we hear singing: "Glory to the Righteous One." But I said, "I waste away, I waste away! Woe to me! The treacherous betray! With treachery the treacherous betray!"
ISA|24|17|Terror and pit and snare await you, O people of the earth.
ISA|24|18|Whoever flees at the sound of terror will fall into a pit; whoever climbs out of the pit will be caught in a snare. The floodgates of the heavens are opened, the foundations of the earth shake.
ISA|24|19|The earth is broken up, the earth is split asunder, the earth is thoroughly shaken.
ISA|24|20|The earth reels like a drunkard, it sways like a hut in the wind; so heavy upon it is the guilt of its rebellion that it falls-never to rise again.
ISA|24|21|In that day the LORD will punish the powers in the heavens above and the kings on the earth below.
ISA|24|22|They will be herded together like prisoners bound in a dungeon; they will be shut up in prison and be punished after many days.
ISA|24|23|The moon will be abashed, the sun ashamed; for the LORD Almighty will reign on Mount Zion and in Jerusalem, and before its elders, gloriously.
ISA|25|1|O LORD, you are my God; I will exalt you and praise your name, for in perfect faithfulness you have done marvelous things, things planned long ago.
ISA|25|2|You have made the city a heap of rubble, the fortified town a ruin, the foreigners' stronghold a city no more; it will never be rebuilt.
ISA|25|3|Therefore strong peoples will honor you; cities of ruthless nations will revere you.
ISA|25|4|You have been a refuge for the poor, a refuge for the needy in his distress, a shelter from the storm and a shade from the heat. For the breath of the ruthless is like a storm driving against a wall
ISA|25|5|and like the heat of the desert. You silence the uproar of foreigners; as heat is reduced by the shadow of a cloud, so the song of the ruthless is stilled.
ISA|25|6|On this mountain the LORD Almighty will prepare a feast of rich food for all peoples, a banquet of aged wine- the best of meats and the finest of wines.
ISA|25|7|On this mountain he will destroy the shroud that enfolds all peoples, the sheet that covers all nations;
ISA|25|8|he will swallow up death forever. The Sovereign LORD will wipe away the tears from all faces; he will remove the disgrace of his people from all the earth. The LORD has spoken.
ISA|25|9|In that day they will say, "Surely this is our God; we trusted in him, and he saved us. This is the LORD, we trusted in him; let us rejoice and be glad in his salvation."
ISA|25|10|The hand of the LORD will rest on this mountain; but Moab will be trampled under him as straw is trampled down in the manure.
ISA|25|11|They will spread out their hands in it, as a swimmer spreads out his hands to swim. God will bring down their pride despite the cleverness of their hands.
ISA|25|12|He will bring down your high fortified walls and lay them low; he will bring them down to the ground, to the very dust.
ISA|26|1|In that day this song will be sung in the land of Judah: We have a strong city; God makes salvation its walls and ramparts.
ISA|26|2|Open the gates that the righteous nation may enter, the nation that keeps faith.
ISA|26|3|You will keep in perfect peace him whose mind is steadfast, because he trusts in you.
ISA|26|4|Trust in the LORD forever, for the LORD, the LORD, is the Rock eternal.
ISA|26|5|He humbles those who dwell on high, he lays the lofty city low; he levels it to the ground and casts it down to the dust.
ISA|26|6|Feet trample it down- the feet of the oppressed, the footsteps of the poor.
ISA|26|7|The path of the righteous is level; O upright One, you make the way of the righteous smooth.
ISA|26|8|Yes, LORD, walking in the way of your laws, we wait for you; your name and renown are the desire of our hearts.
ISA|26|9|My soul yearns for you in the night; in the morning my spirit longs for you. When your judgments come upon the earth, the people of the world learn righteousness.
ISA|26|10|Though grace is shown to the wicked, they do not learn righteousness; even in a land of uprightness they go on doing evil and regard not the majesty of the LORD.
ISA|26|11|O LORD, your hand is lifted high, but they do not see it. Let them see your zeal for your people and be put to shame; let the fire reserved for your enemies consume them.
ISA|26|12|LORD, you establish peace for us; all that we have accomplished you have done for us.
ISA|26|13|O LORD, our God, other lords besides you have ruled over us, but your name alone do we honor.
ISA|26|14|They are now dead, they live no more; those departed spirits do not rise. You punished them and brought them to ruin; you wiped out all memory of them.
ISA|26|15|You have enlarged the nation, O LORD; you have enlarged the nation. You have gained glory for yourself; you have extended all the borders of the land.
ISA|26|16|LORD, they came to you in their distress; when you disciplined them, they could barely whisper a prayer.
ISA|26|17|As a woman with child and about to give birth writhes and cries out in her pain, so were we in your presence, O LORD.
ISA|26|18|We were with child, we writhed in pain, but we gave birth to wind. We have not brought salvation to the earth; we have not given birth to people of the world.
ISA|26|19|But your dead will live; their bodies will rise. You who dwell in the dust, wake up and shout for joy. Your dew is like the dew of the morning; the earth will give birth to her dead.
ISA|26|20|Go, my people, enter your rooms and shut the doors behind you; hide yourselves for a little while until his wrath has passed by.
ISA|26|21|See, the LORD is coming out of his dwelling to punish the people of the earth for their sins. The earth will disclose the blood shed upon her; she will conceal her slain no longer.
ISA|27|1|In that day, the LORD will punish with his sword, his fierce, great and powerful sword, Leviathan the gliding serpent, Leviathan the coiling serpent; he will slay the monster of the sea.
ISA|27|2|In that day- "Sing about a fruitful vineyard:
ISA|27|3|I, the LORD, watch over it; I water it continually. I guard it day and night so that no one may harm it.
ISA|27|4|I am not angry. If only there were briers and thorns confronting me! I would march against them in battle; I would set them all on fire.
ISA|27|5|Or else let them come to me for refuge; let them make peace with me, yes, let them make peace with me."
ISA|27|6|In days to come Jacob will take root, Israel will bud and blossom and fill all the world with fruit.
ISA|27|7|Has the LORD struck her as he struck down those who struck her? Has she been killed as those were killed who killed her?
ISA|27|8|By warfare and exile you contend with her- with his fierce blast he drives her out, as on a day the east wind blows.
ISA|27|9|By this, then, will Jacob's guilt be atoned for, and this will be the full fruitage of the removal of his sin: When he makes all the altar stones to be like chalk stones crushed to pieces, no Asherah poles or incense altars will be left standing.
ISA|27|10|The fortified city stands desolate, an abandoned settlement, forsaken like the desert; there the calves graze, there they lie down; they strip its branches bare.
ISA|27|11|When its twigs are dry, they are broken off and women come and make fires with them. For this is a people without understanding; so their Maker has no compassion on them, and their Creator shows them no favor.
ISA|27|12|In that day the LORD will thresh from the flowing Euphrates to the Wadi of Egypt, and you, O Israelites, will be gathered up one by one.
ISA|27|13|And in that day a great trumpet will sound. Those who were perishing in Assyria and those who were exiled in Egypt will come and worship the LORD on the holy mountain in Jerusalem.
ISA|28|1|Woe to that wreath, the pride of Ephraim's drunkards, to the fading flower, his glorious beauty, set on the head of a fertile valley- to that city, the pride of those laid low by wine!
ISA|28|2|See, the Lord has one who is powerful and strong. Like a hailstorm and a destructive wind, like a driving rain and a flooding downpour, he will throw it forcefully to the ground.
ISA|28|3|That wreath, the pride of Ephraim's drunkards, will be trampled underfoot.
ISA|28|4|That fading flower, his glorious beauty, set on the head of a fertile valley, will be like a fig ripe before harvest- as soon as someone sees it and takes it in his hand, he swallows it.
ISA|28|5|In that day the LORD Almighty will be a glorious crown, a beautiful wreath for the remnant of his people.
ISA|28|6|He will be a spirit of justice to him who sits in judgment, a source of strength to those who turn back the battle at the gate.
ISA|28|7|And these also stagger from wine and reel from beer: Priests and prophets stagger from beer and are befuddled with wine; they reel from beer, they stagger when seeing visions, they stumble when rendering decisions.
ISA|28|8|All the tables are covered with vomit and there is not a spot without filth.
ISA|28|9|"Who is it he is trying to teach? To whom is he explaining his message? To children weaned from their milk, to those just taken from the breast?
ISA|28|10|For it is: Do and do, do and do, rule on rule, rule on rule; a little here, a little there."
ISA|28|11|Very well then, with foreign lips and strange tongues God will speak to this people,
ISA|28|12|to whom he said, "This is the resting place, let the weary rest"; and, "This is the place of repose"- but they would not listen.
ISA|28|13|So then, the word of the LORD to them will become: Do and do, do and do, rule on rule, rule on rule; a little here, a little there- so that they will go and fall backward, be injured and snared and captured.
ISA|28|14|Therefore hear the word of the LORD, you scoffers who rule this people in Jerusalem.
ISA|28|15|You boast, "We have entered into a covenant with death, with the grave we have made an agreement. When an overwhelming scourge sweeps by, it cannot touch us, for we have made a lie our refuge and falsehood our hiding place."
ISA|28|16|So this is what the Sovereign LORD says: "See, I lay a stone in Zion, a tested stone, a precious cornerstone for a sure foundation; the one who trusts will never be dismayed.
ISA|28|17|I will make justice the measuring line and righteousness the plumb line; hail will sweep away your refuge, the lie, and water will overflow your hiding place.
ISA|28|18|Your covenant with death will be annulled; your agreement with the grave will not stand. When the overwhelming scourge sweeps by, you will be beaten down by it.
ISA|28|19|As often as it comes it will carry you away; morning after morning, by day and by night, it will sweep through." The understanding of this message will bring sheer terror.
ISA|28|20|The bed is too short to stretch out on, the blanket too narrow to wrap around you.
ISA|28|21|The LORD will rise up as he did at Mount Perazim, he will rouse himself as in the Valley of Gibeon- to do his work, his strange work, and perform his task, his alien task.
ISA|28|22|Now stop your mocking, or your chains will become heavier; the Lord, the LORD Almighty, has told me of the destruction decreed against the whole land.
ISA|28|23|Listen and hear my voice; pay attention and hear what I say.
ISA|28|24|When a farmer plows for planting, does he plow continually? Does he keep on breaking up and harrowing the soil?
ISA|28|25|When he has leveled the surface, does he not sow caraway and scatter cummin? Does he not plant wheat in its place, barley in its plot, and spelt in its field?
ISA|28|26|His God instructs him and teaches him the right way.
ISA|28|27|Caraway is not threshed with a sledge, nor is a cartwheel rolled over cummin; caraway is beaten out with a rod, and cummin with a stick.
ISA|28|28|Grain must be ground to make bread; so one does not go on threshing it forever. Though he drives the wheels of his threshing cart over it, his horses do not grind it.
ISA|28|29|All this also comes from the LORD Almighty, wonderful in counsel and magnificent in wisdom.
ISA|29|1|Woe to you, Ariel, Ariel, the city where David settled! Add year to year and let your cycle of festivals go on.
ISA|29|2|Yet I will besiege Ariel; she will mourn and lament, she will be to me like an altar hearth.
ISA|29|3|I will encamp against you all around; I will encircle you with towers and set up my siege works against you.
ISA|29|4|Brought low, you will speak from the ground; your speech will mumble out of the dust. Your voice will come ghostlike from the earth; out of the dust your speech will whisper.
ISA|29|5|But your many enemies will become like fine dust, the ruthless hordes like blown chaff. Suddenly, in an instant,
ISA|29|6|the LORD Almighty will come with thunder and earthquake and great noise, with windstorm and tempest and flames of a devouring fire.
ISA|29|7|Then the hordes of all the nations that fight against Ariel, that attack her and her fortress and besiege her, will be as it is with a dream, with a vision in the night-
ISA|29|8|as when a hungry man dreams that he is eating, but he awakens, and his hunger remains; as when a thirsty man dreams that he is drinking, but he awakens faint, with his thirst unquenched. So will it be with the hordes of all the nations that fight against Mount Zion.
ISA|29|9|Be stunned and amazed, blind yourselves and be sightless; be drunk, but not from wine, stagger, but not from beer.
ISA|29|10|The LORD has brought over you a deep sleep: He has sealed your eyes (the prophets); he has covered your heads (the seers).
ISA|29|11|For you this whole vision is nothing but words sealed in a scroll. And if you give the scroll to someone who can read, and say to him, "Read this, please," he will answer, "I can't; it is sealed."
ISA|29|12|Or if you give the scroll to someone who cannot read, and say, "Read this, please," he will answer, "I don't know how to read."
ISA|29|13|The Lord says: "These people come near to me with their mouth and honor me with their lips, but their hearts are far from me. Their worship of me is made up only of rules taught by men.
ISA|29|14|Therefore once more I will astound these people with wonder upon wonder; the wisdom of the wise will perish, the intelligence of the intelligent will vanish."
ISA|29|15|Woe to those who go to great depths to hide their plans from the LORD, who do their work in darkness and think, "Who sees us? Who will know?"
ISA|29|16|You turn things upside down, as if the potter were thought to be like the clay! Shall what is formed say to him who formed it, "He did not make me"? Can the pot say of the potter, "He knows nothing"?
ISA|29|17|In a very short time, will not Lebanon be turned into a fertile field and the fertile field seem like a forest?
ISA|29|18|In that day the deaf will hear the words of the scroll, and out of gloom and darkness the eyes of the blind will see.
ISA|29|19|Once more the humble will rejoice in the LORD; the needy will rejoice in the Holy One of Israel.
ISA|29|20|The ruthless will vanish, the mockers will disappear, and all who have an eye for evil will be cut down-
ISA|29|21|those who with a word make a man out to be guilty, who ensnare the defender in court and with false testimony deprive the innocent of justice.
ISA|29|22|Therefore this is what the LORD, who redeemed Abraham, says to the house of Jacob: "No longer will Jacob be ashamed; no longer will their faces grow pale.
ISA|29|23|When they see among them their children, the work of my hands, they will keep my name holy; they will acknowledge the holiness of the Holy One of Jacob, and will stand in awe of the God of Israel.
ISA|29|24|Those who are wayward in spirit will gain understanding; those who complain will accept instruction."
ISA|30|1|"Woe to the obstinate children," declares the LORD, "to those who carry out plans that are not mine, forming an alliance, but not by my Spirit, heaping sin upon sin;
ISA|30|2|who go down to Egypt without consulting me; who look for help to Pharaoh's protection, to Egypt's shade for refuge.
ISA|30|3|But Pharaoh's protection will be to your shame, Egypt's shade will bring you disgrace.
ISA|30|4|Though they have officials in Zoan and their envoys have arrived in Hanes,
ISA|30|5|everyone will be put to shame because of a people useless to them, who bring neither help nor advantage, but only shame and disgrace."
ISA|30|6|An oracle concerning the animals of the Negev: Through a land of hardship and distress, of lions and lionesses, of adders and darting snakes, the envoys carry their riches on donkeys' backs, their treasures on the humps of camels, to that unprofitable nation,
ISA|30|7|to Egypt, whose help is utterly useless. Therefore I call her Rahab the Do-Nothing.
ISA|30|8|Go now, write it on a tablet for them, inscribe it on a scroll, that for the days to come it may be an everlasting witness.
ISA|30|9|These are rebellious people, deceitful children, children unwilling to listen to the LORD's instruction.
ISA|30|10|They say to the seers, "See no more visions!" and to the prophets, "Give us no more visions of what is right! Tell us pleasant things, prophesy illusions.
ISA|30|11|Leave this way, get off this path, and stop confronting us with the Holy One of Israel!"
ISA|30|12|Therefore, this is what the Holy One of Israel says: "Because you have rejected this message, relied on oppression and depended on deceit,
ISA|30|13|this sin will become for you like a high wall, cracked and bulging, that collapses suddenly, in an instant.
ISA|30|14|It will break in pieces like pottery, shattered so mercilessly that among its pieces not a fragment will be found for taking coals from a hearth or scooping water out of a cistern."
ISA|30|15|This is what the Sovereign LORD, the Holy One of Israel, says: "In repentance and rest is your salvation, in quietness and trust is your strength, but you would have none of it.
ISA|30|16|You said, 'No, we will flee on horses.' Therefore you will flee! You said, 'We will ride off on swift horses.' Therefore your pursuers will be swift!
ISA|30|17|A thousand will flee at the threat of one; at the threat of five you will all flee away, till you are left like a flagstaff on a mountaintop, like a banner on a hill."
ISA|30|18|Yet the LORD longs to be gracious to you; he rises to show you compassion. For the LORD is a God of justice. Blessed are all who wait for him!
ISA|30|19|O people of Zion, who live in Jerusalem, you will weep no more. How gracious he will be when you cry for help! As soon as he hears, he will answer you.
ISA|30|20|Although the Lord gives you the bread of adversity and the water of affliction, your teachers will be hidden no more; with your own eyes you will see them.
ISA|30|21|Whether you turn to the right or to the left, your ears will hear a voice behind you, saying, "This is the way; walk in it."
ISA|30|22|Then you will defile your idols overlaid with silver and your images covered with gold; you will throw them away like a menstrual cloth and say to them, "Away with you!"
ISA|30|23|He will also send you rain for the seed you sow in the ground, and the food that comes from the land will be rich and plentiful. In that day your cattle will graze in broad meadows.
ISA|30|24|The oxen and donkeys that work the soil will eat fodder and mash, spread out with fork and shovel.
ISA|30|25|In the day of great slaughter, when the towers fall, streams of water will flow on every high mountain and every lofty hill.
ISA|30|26|The moon will shine like the sun, and the sunlight will be seven times brighter, like the light of seven full days, when the LORD binds up the bruises of his people and heals the wounds he inflicted.
ISA|30|27|See, the Name of the LORD comes from afar, with burning anger and dense clouds of smoke; his lips are full of wrath, and his tongue is a consuming fire.
ISA|30|28|His breath is like a rushing torrent, rising up to the neck. He shakes the nations in the sieve of destruction; he places in the jaws of the peoples a bit that leads them astray.
ISA|30|29|And you will sing as on the night you celebrate a holy festival; your hearts will rejoice as when people go up with flutes to the mountain of the LORD, to the Rock of Israel.
ISA|30|30|The LORD will cause men to hear his majestic voice and will make them see his arm coming down with raging anger and consuming fire, with cloudburst, thunderstorm and hail.
ISA|30|31|The voice of the LORD will shatter Assyria; with his scepter he will strike them down.
ISA|30|32|Every stroke the LORD lays on them with his punishing rod will be to the music of tambourines and harps, as he fights them in battle with the blows of his arm.
ISA|30|33|Topheth has long been prepared; it has been made ready for the king. Its fire pit has been made deep and wide, with an abundance of fire and wood; the breath of the LORD, like a stream of burning sulfur, sets it ablaze.
ISA|31|1|Woe to those who go down to Egypt for help, who rely on horses, who trust in the multitude of their chariots and in the great strength of their horsemen, but do not look to the Holy One of Israel, or seek help from the LORD.
ISA|31|2|Yet he too is wise and can bring disaster; he does not take back his words. He will rise up against the house of the wicked, against those who help evildoers.
ISA|31|3|But the Egyptians are men and not God; their horses are flesh and not spirit. When the LORD stretches out his hand, he who helps will stumble, he who is helped will fall; both will perish together.
ISA|31|4|This is what the LORD says to me: "As a lion growls, a great lion over his prey- and though a whole band of shepherds is called together against him, he is not frightened by their shouts or disturbed by their clamor- so the LORD Almighty will come down to do battle on Mount Zion and on its heights.
ISA|31|5|Like birds hovering overhead, the LORD Almighty will shield Jerusalem; he will shield it and deliver it, he will 'pass over' it and will rescue it."
ISA|31|6|Return to him you have so greatly revolted against, O Israelites.
ISA|31|7|For in that day every one of you will reject the idols of silver and gold your sinful hands have made.
ISA|31|8|"Assyria will fall by a sword that is not of man; a sword, not of mortals, will devour them. They will flee before the sword and their young men will be put to forced labor.
ISA|31|9|Their stronghold will fall because of terror; at sight of the battle standard their commanders will panic," declares the LORD, whose fire is in Zion, whose furnace is in Jerusalem.
ISA|32|1|See, a king will reign in righteousness and rulers will rule with justice.
ISA|32|2|Each man will be like a shelter from the wind and a refuge from the storm, like streams of water in the desert and the shadow of a great rock in a thirsty land.
ISA|32|3|Then the eyes of those who see will no longer be closed, and the ears of those who hear will listen.
ISA|32|4|The mind of the rash will know and understand, and the stammering tongue will be fluent and clear.
ISA|32|5|No longer will the fool be called noble nor the scoundrel be highly respected.
ISA|32|6|For the fool speaks folly, his mind is busy with evil: He practices ungodliness and spreads error concerning the LORD; the hungry he leaves empty and from the thirsty he withholds water.
ISA|32|7|The scoundrel's methods are wicked, he makes up evil schemes to destroy the poor with lies, even when the plea of the needy is just.
ISA|32|8|But the noble man makes noble plans, and by noble deeds he stands.
ISA|32|9|You women who are so complacent, rise up and listen to me; you daughters who feel secure, hear what I have to say!
ISA|32|10|In little more than a year you who feel secure will tremble; the grape harvest will fail, and the harvest of fruit will not come.
ISA|32|11|Tremble, you complacent women; shudder, you daughters who feel secure! Strip off your clothes, put sackcloth around your waists.
ISA|32|12|Beat your breasts for the pleasant fields, for the fruitful vines
ISA|32|13|and for the land of my people, a land overgrown with thorns and briers- yes, mourn for all houses of merriment and for this city of revelry.
ISA|32|14|The fortress will be abandoned, the noisy city deserted; citadel and watchtower will become a wasteland forever, the delight of donkeys, a pasture for flocks,
ISA|32|15|till the Spirit is poured upon us from on high, and the desert becomes a fertile field, and the fertile field seems like a forest.
ISA|32|16|Justice will dwell in the desert and righteousness live in the fertile field.
ISA|32|17|The fruit of righteousness will be peace; the effect of righteousness will be quietness and confidence forever.
ISA|32|18|My people will live in peaceful dwelling places, in secure homes, in undisturbed places of rest.
ISA|32|19|Though hail flattens the forest and the city is leveled completely,
ISA|32|20|how blessed you will be, sowing your seed by every stream, and letting your cattle and donkeys range free.
ISA|33|1|Woe to you, O destroyer, you who have not been destroyed! Woe to you, O traitor, you who have not been betrayed! When you stop destroying, you will be destroyed; when you stop betraying, you will be betrayed.
ISA|33|2|O LORD, be gracious to us; we long for you. Be our strength every morning, our salvation in time of distress.
ISA|33|3|At the thunder of your voice, the peoples flee; when you rise up, the nations scatter.
ISA|33|4|Your plunder, O nations, is harvested as by young locusts; like a swarm of locusts men pounce on it.
ISA|33|5|The LORD is exalted, for he dwells on high; he will fill Zion with justice and righteousness.
ISA|33|6|He will be the sure foundation for your times, a rich store of salvation and wisdom and knowledge; the fear of the LORD is the key to this treasure.
ISA|33|7|Look, their brave men cry aloud in the streets; the envoys of peace weep bitterly.
ISA|33|8|The highways are deserted, no travelers are on the roads. The treaty is broken, its witnesses are despised, no one is respected.
ISA|33|9|The land mourns and wastes away, Lebanon is ashamed and withers; Sharon is like the Arabah, and Bashan and Carmel drop their leaves.
ISA|33|10|"Now will I arise," says the LORD. "Now will I be exalted; now will I be lifted up.
ISA|33|11|You conceive chaff, you give birth to straw; your breath is a fire that consumes you.
ISA|33|12|The peoples will be burned as if to lime; like cut thornbushes they will be set ablaze."
ISA|33|13|You who are far away, hear what I have done; you who are near, acknowledge my power!
ISA|33|14|The sinners in Zion are terrified; trembling grips the godless: "Who of us can dwell with the consuming fire? Who of us can dwell with everlasting burning?"
ISA|33|15|He who walks righteously and speaks what is right, who rejects gain from extortion and keeps his hand from accepting bribes, who stops his ears against plots of murder and shuts his eyes against contemplating evil-
ISA|33|16|this is the man who will dwell on the heights, whose refuge will be the mountain fortress. His bread will be supplied, and water will not fail him.
ISA|33|17|Your eyes will see the king in his beauty and view a land that stretches afar.
ISA|33|18|In your thoughts you will ponder the former terror: "Where is that chief officer? Where is the one who took the revenue? Where is the officer in charge of the towers?"
ISA|33|19|You will see those arrogant people no more, those people of an obscure speech, with their strange, incomprehensible tongue.
ISA|33|20|Look upon Zion, the city of our festivals; your eyes will see Jerusalem, a peaceful abode, a tent that will not be moved; its stakes will never be pulled up, nor any of its ropes broken.
ISA|33|21|There the LORD will be our Mighty One. It will be like a place of broad rivers and streams. No galley with oars will ride them, no mighty ship will sail them.
ISA|33|22|For the LORD is our judge, the LORD is our lawgiver, the LORD is our king; it is he who will save us.
ISA|33|23|Your rigging hangs loose: The mast is not held secure, the sail is not spread. Then an abundance of spoils will be divided and even the lame will carry off plunder.
ISA|33|24|No one living in Zion will say, "I am ill"; and the sins of those who dwell there will be forgiven.
ISA|34|1|Come near, you nations, and listen; pay attention, you peoples! Let the earth hear, and all that is in it, the world, and all that comes out of it!
ISA|34|2|The LORD is angry with all nations; his wrath is upon all their armies. He will totally destroy them, he will give them over to slaughter.
ISA|34|3|Their slain will be thrown out, their dead bodies will send up a stench; the mountains will be soaked with their blood.
ISA|34|4|All the stars of the heavens will be dissolved and the sky rolled up like a scroll; all the starry host will fall like withered leaves from the vine, like shriveled figs from the fig tree.
ISA|34|5|My sword has drunk its fill in the heavens; see, it descends in judgment on Edom, the people I have totally destroyed.
ISA|34|6|The sword of the LORD is bathed in blood, it is covered with fat- the blood of lambs and goats, fat from the kidneys of rams. For the LORD has a sacrifice in Bozrah and a great slaughter in Edom.
ISA|34|7|And the wild oxen will fall with them, the bull calves and the great bulls. Their land will be drenched with blood, and the dust will be soaked with fat.
ISA|34|8|For the LORD has a day of vengeance, a year of retribution, to uphold Zion's cause.
ISA|34|9|Edom's streams will be turned into pitch, her dust into burning sulfur; her land will become blazing pitch!
ISA|34|10|It will not be quenched night and day; its smoke will rise forever. From generation to generation it will lie desolate; no one will ever pass through it again.
ISA|34|11|The desert owl and screech owl will possess it; the great owl and the raven will nest there. God will stretch out over Edom the measuring line of chaos and the plumb line of desolation.
ISA|34|12|Her nobles will have nothing there to be called a kingdom, all her princes will vanish away.
ISA|34|13|Thorns will overrun her citadels, nettles and brambles her strongholds. She will become a haunt for jackals, a home for owls.
ISA|34|14|Desert creatures will meet with hyenas, and wild goats will bleat to each other; there the night creatures will also repose and find for themselves places of rest.
ISA|34|15|The owl will nest there and lay eggs, she will hatch them, and care for her young under the shadow of her wings; there also the falcons will gather, each with its mate.
ISA|34|16|Look in the scroll of the LORD and read: None of these will be missing, not one will lack her mate. For it is his mouth that has given the order, and his Spirit will gather them together.
ISA|34|17|He allots their portions; his hand distributes them by measure. They will possess it forever and dwell there from generation to generation.
ISA|35|1|The desert and the parched land will be glad; the wilderness will rejoice and blossom. Like the crocus,
ISA|35|2|it will burst into bloom; it will rejoice greatly and shout for joy. The glory of Lebanon will be given to it, the splendor of Carmel and Sharon; they will see the glory of the LORD, the splendor of our God.
ISA|35|3|Strengthen the feeble hands, steady the knees that give way;
ISA|35|4|say to those with fearful hearts, "Be strong, do not fear; your God will come, he will come with vengeance; with divine retribution he will come to save you."
ISA|35|5|Then will the eyes of the blind be opened and the ears of the deaf unstopped.
ISA|35|6|Then will the lame leap like a deer, and the mute tongue shout for joy. Water will gush forth in the wilderness and streams in the desert.
ISA|35|7|The burning sand will become a pool, the thirsty ground bubbling springs. In the haunts where jackals once lay, grass and reeds and papyrus will grow.
ISA|35|8|And a highway will be there; it will be called the Way of Holiness. The unclean will not journey on it; it will be for those who walk in that Way; wicked fools will not go about on it.
ISA|35|9|No lion will be there, nor will any ferocious beast get up on it; they will not be found there. But only the redeemed will walk there,
ISA|35|10|and the ransomed of the LORD will return. They will enter Zion with singing; everlasting joy will crown their heads. Gladness and joy will overtake them, and sorrow and sighing will flee away.
ISA|36|1|In the fourteenth year of King Hezekiah's reign, Sennacherib king of Assyria attacked all the fortified cities of Judah and captured them.
ISA|36|2|Then the king of Assyria sent his field commander with a large army from Lachish to King Hezekiah at Jerusalem. When the commander stopped at the aqueduct of the Upper Pool, on the road to the Washerman's Field,
ISA|36|3|Eliakim son of Hilkiah the palace administrator, Shebna the secretary, and Joah son of Asaph the recorder went out to him.
ISA|36|4|The field commander said to them, "Tell Hezekiah, "'This is what the great king, the king of Assyria, says: On what are you basing this confidence of yours?
ISA|36|5|You say you have strategy and military strength-but you speak only empty words. On whom are you depending, that you rebel against me?
ISA|36|6|Look now, you are depending on Egypt, that splintered reed of a staff, which pierces a man's hand and wounds him if he leans on it! Such is Pharaoh king of Egypt to all who depend on him.
ISA|36|7|And if you say to me, "We are depending on the LORD our God"-isn't he the one whose high places and altars Hezekiah removed, saying to Judah and Jerusalem, "You must worship before this altar"?
ISA|36|8|"'Come now, make a bargain with my master, the king of Assyria: I will give you two thousand horses-if you can put riders on them!
ISA|36|9|How then can you repulse one officer of the least of my master's officials, even though you are depending on Egypt for chariots and horsemen?
ISA|36|10|Furthermore, have I come to attack and destroy this land without the LORD? The LORD himself told me to march against this country and destroy it.'"
ISA|36|11|Then Eliakim, Shebna and Joah said to the field commander, "Please speak to your servants in Aramaic, since we understand it. Don't speak to us in Hebrew in the hearing of the people on the wall."
ISA|36|12|But the commander replied, "Was it only to your master and you that my master sent me to say these things, and not to the men sitting on the wall-who, like you, will have to eat their own filth and drink their own urine?"
ISA|36|13|Then the commander stood and called out in Hebrew, "Hear the words of the great king, the king of Assyria!
ISA|36|14|This is what the king says: Do not let Hezekiah deceive you. He cannot deliver you!
ISA|36|15|Do not let Hezekiah persuade you to trust in the LORD when he says, 'The LORD will surely deliver us; this city will not be given into the hand of the king of Assyria.'
ISA|36|16|"Do not listen to Hezekiah. This is what the king of Assyria says: Make peace with me and come out to me. Then every one of you will eat from his own vine and fig tree and drink water from his own cistern,
ISA|36|17|until I come and take you to a land like your own-a land of grain and new wine, a land of bread and vineyards.
ISA|36|18|"Do not let Hezekiah mislead you when he says, 'The LORD will deliver us.' Has the god of any nation ever delivered his land from the hand of the king of Assyria?
ISA|36|19|Where are the gods of Hamath and Arpad? Where are the gods of Sepharvaim? Have they rescued Samaria from my hand?
ISA|36|20|Who of all the gods of these countries has been able to save his land from me? How then can the LORD deliver Jerusalem from my hand?"
ISA|36|21|But the people remained silent and said nothing in reply, because the king had commanded, "Do not answer him."
ISA|36|22|Then Eliakim son of Hilkiah the palace administrator, Shebna the secretary, and Joah son of Asaph the recorder went to Hezekiah, with their clothes torn, and told him what the field commander had said.
ISA|37|1|When King Hezekiah heard this, he tore his clothes and put on sackcloth and went into the temple of the LORD.
ISA|37|2|He sent Eliakim the palace administrator, Shebna the secretary, and the leading priests, all wearing sackcloth, to the prophet Isaiah son of Amoz.
ISA|37|3|They told him, "This is what Hezekiah says: This day is a day of distress and rebuke and disgrace, as when children come to the point of birth and there is no strength to deliver them.
ISA|37|4|It may be that the LORD your God will hear the words of the field commander, whom his master, the king of Assyria, has sent to ridicule the living God, and that he will rebuke him for the words the LORD your God has heard. Therefore pray for the remnant that still survives."
ISA|37|5|When King Hezekiah's officials came to Isaiah,
ISA|37|6|Isaiah said to them, "Tell your master, 'This is what the LORD says: Do not be afraid of what you have heard-those words with which the underlings of the king of Assyria have blasphemed me.
ISA|37|7|Listen! I am going to put a spirit in him so that when he hears a certain report, he will return to his own country, and there I will have him cut down with the sword.'"
ISA|37|8|When the field commander heard that the king of Assyria had left Lachish, he withdrew and found the king fighting against Libnah.
ISA|37|9|Now Sennacherib received a report that Tirhakah, the Cushite king of Egypt, was marching out to fight against him. When he heard it, he sent messengers to Hezekiah with this word:
ISA|37|10|"Say to Hezekiah king of Judah: Do not let the god you depend on deceive you when he says, 'Jerusalem will not be handed over to the king of Assyria.'
ISA|37|11|Surely you have heard what the kings of Assyria have done to all the countries, destroying them completely. And will you be delivered?
ISA|37|12|Did the gods of the nations that were destroyed by my forefathers deliver them-the gods of Gozan, Haran, Rezeph and the people of Eden who were in Tel Assar?
ISA|37|13|Where is the king of Hamath, the king of Arpad, the king of the city of Sepharvaim, or of Hena or Ivvah?"
ISA|37|14|Hezekiah received the letter from the messengers and read it. Then he went up to the temple of the LORD and spread it out before the LORD.
ISA|37|15|And Hezekiah prayed to the LORD:
ISA|37|16|"O LORD Almighty, God of Israel, enthroned between the cherubim, you alone are God over all the kingdoms of the earth. You have made heaven and earth.
ISA|37|17|Give ear, O LORD, and hear; open your eyes, O LORD, and see; listen to all the words Sennacherib has sent to insult the living God.
ISA|37|18|"It is true, O LORD, that the Assyrian kings have laid waste all these peoples and their lands.
ISA|37|19|They have thrown their gods into the fire and destroyed them, for they were not gods but only wood and stone, fashioned by human hands.
ISA|37|20|Now, O LORD our God, deliver us from his hand, so that all kingdoms on earth may know that you alone, O LORD, are God. "
ISA|37|21|Then Isaiah son of Amoz sent a message to Hezekiah: "This is what the LORD, the God of Israel, says: Because you have prayed to me concerning Sennacherib king of Assyria,
ISA|37|22|this is the word the LORD has spoken against him: "The Virgin Daughter of Zion despises and mocks you. The Daughter of Jerusalem tosses her head as you flee.
ISA|37|23|Who is it you have insulted and blasphemed? Against whom have you raised your voice and lifted your eyes in pride? Against the Holy One of Israel!
ISA|37|24|By your messengers you have heaped insults on the Lord. And you have said, 'With my many chariots I have ascended the heights of the mountains, the utmost heights of Lebanon. I have cut down its tallest cedars, the choicest of its pines. I have reached its remotest heights, the finest of its forests.
ISA|37|25|I have dug wells in foreign lands and drunk the water there. With the soles of my feet I have dried up all the streams of Egypt.'
ISA|37|26|"Have you not heard? Long ago I ordained it. In days of old I planned it; now I have brought it to pass, that you have turned fortified cities into piles of stone.
ISA|37|27|Their people, drained of power, are dismayed and put to shame. They are like plants in the field, like tender green shoots, like grass sprouting on the roof, scorched before it grows up.
ISA|37|28|"But I know where you stay and when you come and go and how you rage against me.
ISA|37|29|Because you rage against me and because your insolence has reached my ears, I will put my hook in your nose and my bit in your mouth, and I will make you return by the way you came.
ISA|37|30|"This will be the sign for you, O Hezekiah: "This year you will eat what grows by itself, and the second year what springs from that. But in the third year sow and reap, plant vineyards and eat their fruit.
ISA|37|31|Once more a remnant of the house of Judah will take root below and bear fruit above.
ISA|37|32|For out of Jerusalem will come a remnant, and out of Mount Zion a band of survivors. The zeal of the LORD Almighty will accomplish this.
ISA|37|33|"Therefore this is what the LORD says concerning the king of Assyria: "He will not enter this city or shoot an arrow here. He will not come before it with shield or build a siege ramp against it.
ISA|37|34|By the way that he came he will return; he will not enter this city," declares the LORD.
ISA|37|35|"I will defend this city and save it, for my sake and for the sake of David my servant!"
ISA|37|36|Then the angel of the LORD went out and put to death a hundred and eighty-five thousand men in the Assyrian camp. When the people got up the next morning-there were all the dead bodies!
ISA|37|37|So Sennacherib king of Assyria broke camp and withdrew. He returned to Nineveh and stayed there.
ISA|37|38|One day, while he was worshiping in the temple of his god Nisroch, his sons Adrammelech and Sharezer cut him down with the sword, and they escaped to the land of Ararat. And Esarhaddon his son succeeded him as king.
ISA|38|1|In those days Hezekiah became ill and was at the point of death. The prophet Isaiah son of Amoz went to him and said, "This is what the LORD says: Put your house in order, because you are going to die; you will not recover."
ISA|38|2|Hezekiah turned his face to the wall and prayed to the LORD,
ISA|38|3|"Remember, O LORD, how I have walked before you faithfully and with wholehearted devotion and have done what is good in your eyes." And Hezekiah wept bitterly.
ISA|38|4|Then the word of the LORD came to Isaiah:
ISA|38|5|"Go and tell Hezekiah, 'This is what the LORD, the God of your father David, says: I have heard your prayer and seen your tears; I will add fifteen years to your life.
ISA|38|6|And I will deliver you and this city from the hand of the king of Assyria. I will defend this city.
ISA|38|7|"'This is the LORD's sign to you that the LORD will do what he has promised:
ISA|38|8|I will make the shadow cast by the sun go back the ten steps it has gone down on the stairway of Ahaz.'" So the sunlight went back the ten steps it had gone down.
ISA|38|9|A writing of Hezekiah king of Judah after his illness and recovery:
ISA|38|10|I said, "In the prime of my life must I go through the gates of death and be robbed of the rest of my years?"
ISA|38|11|I said, "I will not again see the LORD, the LORD, in the land of the living; no longer will I look on mankind, or be with those who now dwell in this world.
ISA|38|12|Like a shepherd's tent my house has been pulled down and taken from me. Like a weaver I have rolled up my life, and he has cut me off from the loom; day and night you made an end of me.
ISA|38|13|I waited patiently till dawn, but like a lion he broke all my bones; day and night you made an end of me.
ISA|38|14|I cried like a swift or thrush, I moaned like a mourning dove. My eyes grew weak as I looked to the heavens. I am troubled; O Lord, come to my aid!"
ISA|38|15|But what can I say? He has spoken to me, and he himself has done this. I will walk humbly all my years because of this anguish of my soul.
ISA|38|16|Lord, by such things men live; and my spirit finds life in them too. You restored me to health and let me live.
ISA|38|17|Surely it was for my benefit that I suffered such anguish. In your love you kept me from the pit of destruction; you have put all my sins behind your back.
ISA|38|18|For the grave cannot praise you, death cannot sing your praise; those who go down to the pit cannot hope for your faithfulness.
ISA|38|19|The living, the living-they praise you, as I am doing today; fathers tell their children about your faithfulness.
ISA|38|20|The LORD will save me, and we will sing with stringed instruments all the days of our lives in the temple of the LORD.
ISA|38|21|Isaiah had said, "Prepare a poultice of figs and apply it to the boil, and he will recover."
ISA|38|22|Hezekiah had asked, "What will be the sign that I will go up to the temple of the LORD?"
ISA|39|1|At that time Merodach-Baladan son of Baladan king of Babylon sent Hezekiah letters and a gift, because he had heard of his illness and recovery.
ISA|39|2|Hezekiah received the envoys gladly and showed them what was in his storehouses-the silver, the gold, the spices, the fine oil, his entire armory and everything found among his treasures. There was nothing in his palace or in all his kingdom that Hezekiah did not show them.
ISA|39|3|Then Isaiah the prophet went to King Hezekiah and asked, "What did those men say, and where did they come from?From a distant land," Hezekiah replied. "They came to me from Babylon."
ISA|39|4|The prophet asked, "What did they see in your palace?They saw everything in my palace," Hezekiah said. "There is nothing among my treasures that I did not show them."
ISA|39|5|Then Isaiah said to Hezekiah, "Hear the word of the LORD Almighty:
ISA|39|6|The time will surely come when everything in your palace, and all that your fathers have stored up until this day, will be carried off to Babylon. Nothing will be left, says the LORD.
ISA|39|7|And some of your descendants, your own flesh and blood who will be born to you, will be taken away, and they will become eunuchs in the palace of the king of Babylon."
ISA|39|8|"The word of the LORD you have spoken is good," Hezekiah replied. For he thought, "There will be peace and security in my lifetime."
ISA|40|1|Comfort, comfort my people, says your God.
ISA|40|2|Speak tenderly to Jerusalem, and proclaim to her that her hard service has been completed, that her sin has been paid for, that she has received from the LORD's hand double for all her sins.
ISA|40|3|A voice of one calling: "In the desert prepare the way for the LORD; make straight in the wilderness a highway for our God.
ISA|40|4|Every valley shall be raised up, every mountain and hill made low; the rough ground shall become level, the rugged places a plain.
ISA|40|5|And the glory of the LORD will be revealed, and all mankind together will see it. For the mouth of the LORD has spoken."
ISA|40|6|A voice says, "Cry out." And I said, "What shall I cry?All men are like grass, and all their glory is like the flowers of the field.
ISA|40|7|The grass withers and the flowers fall, because the breath of the LORD blows on them. Surely the people are grass.
ISA|40|8|The grass withers and the flowers fall, but the word of our God stands forever."
ISA|40|9|You who bring good tidings to Zion, go up on a high mountain. You who bring good tidings to Jerusalem, lift up your voice with a shout, lift it up, do not be afraid; say to the towns of Judah, "Here is your God!"
ISA|40|10|See, the Sovereign LORD comes with power, and his arm rules for him. See, his reward is with him, and his recompense accompanies him.
ISA|40|11|He tends his flock like a shepherd: He gathers the lambs in his arms and carries them close to his heart; he gently leads those that have young.
ISA|40|12|Who has measured the waters in the hollow of his hand, or with the breadth of his hand marked off the heavens? Who has held the dust of the earth in a basket, or weighed the mountains on the scales and the hills in a balance?
ISA|40|13|Who has understood the mind of the LORD, or instructed him as his counselor?
ISA|40|14|Whom did the LORD consult to enlighten him, and who taught him the right way? Who was it that taught him knowledge or showed him the path of understanding?
ISA|40|15|Surely the nations are like a drop in a bucket; they are regarded as dust on the scales; he weighs the islands as though they were fine dust.
ISA|40|16|Lebanon is not sufficient for altar fires, nor its animals enough for burnt offerings.
ISA|40|17|Before him all the nations are as nothing; they are regarded by him as worthless and less than nothing.
ISA|40|18|To whom, then, will you compare God? What image will you compare him to?
ISA|40|19|As for an idol, a craftsman casts it, and a goldsmith overlays it with gold and fashions silver chains for it.
ISA|40|20|A man too poor to present such an offering selects wood that will not rot. He looks for a skilled craftsman to set up an idol that will not topple.
ISA|40|21|Do you not know? Have you not heard? Has it not been told you from the beginning? Have you not understood since the earth was founded?
ISA|40|22|He sits enthroned above the circle of the earth, and its people are like grasshoppers. He stretches out the heavens like a canopy, and spreads them out like a tent to live in.
ISA|40|23|He brings princes to naught and reduces the rulers of this world to nothing.
ISA|40|24|No sooner are they planted, no sooner are they sown, no sooner do they take root in the ground, than he blows on them and they wither, and a whirlwind sweeps them away like chaff.
ISA|40|25|"To whom will you compare me? Or who is my equal?" says the Holy One.
ISA|40|26|Lift your eyes and look to the heavens: Who created all these? He who brings out the starry host one by one, and calls them each by name. Because of his great power and mighty strength, not one of them is missing.
ISA|40|27|Why do you say, O Jacob, and complain, O Israel, "My way is hidden from the LORD; my cause is disregarded by my God"?
ISA|40|28|Do you not know? Have you not heard? The LORD is the everlasting God, the Creator of the ends of the earth. He will not grow tired or weary, and his understanding no one can fathom.
ISA|40|29|He gives strength to the weary and increases the power of the weak.
ISA|40|30|Even youths grow tired and weary, and young men stumble and fall;
ISA|40|31|but those who hope in the LORD will renew their strength. They will soar on wings like eagles; they will run and not grow weary, they will walk and not be faint.
ISA|41|1|"Be silent before me, you islands! Let the nations renew their strength! Let them come forward and speak; let us meet together at the place of judgment.
ISA|41|2|"Who has stirred up one from the east, calling him in righteousness to his service? He hands nations over to him and subdues kings before him. He turns them to dust with his sword, to windblown chaff with his bow.
ISA|41|3|He pursues them and moves on unscathed, by a path his feet have not traveled before.
ISA|41|4|Who has done this and carried it through, calling forth the generations from the beginning? I, the LORD -with the first of them and with the last-I am he."
ISA|41|5|The islands have seen it and fear; the ends of the earth tremble. They approach and come forward;
ISA|41|6|each helps the other and says to his brother, "Be strong!"
ISA|41|7|The craftsman encourages the goldsmith, and he who smooths with the hammer spurs on him who strikes the anvil. He says of the welding, "It is good." He nails down the idol so it will not topple.
ISA|41|8|"But you, O Israel, my servant, Jacob, whom I have chosen, you descendants of Abraham my friend,
ISA|41|9|I took you from the ends of the earth, from its farthest corners I called you. I said, 'You are my servant'; I have chosen you and have not rejected you.
ISA|41|10|So do not fear, for I am with you; do not be dismayed, for I am your God. I will strengthen you and help you; I will uphold you with my righteous right hand.
ISA|41|11|"All who rage against you will surely be ashamed and disgraced; those who oppose you will be as nothing and perish.
ISA|41|12|Though you search for your enemies, you will not find them. Those who wage war against you will be as nothing at all.
ISA|41|13|For I am the LORD, your God, who takes hold of your right hand and says to you, Do not fear; I will help you.
ISA|41|14|Do not be afraid, O worm Jacob, O little Israel, for I myself will help you," declares the LORD, your Redeemer, the Holy One of Israel.
ISA|41|15|"See, I will make you into a threshing sledge, new and sharp, with many teeth. You will thresh the mountains and crush them, and reduce the hills to chaff.
ISA|41|16|You will winnow them, the wind will pick them up, and a gale will blow them away. But you will rejoice in the LORD and glory in the Holy One of Israel.
ISA|41|17|"The poor and needy search for water, but there is none; their tongues are parched with thirst. But I the LORD will answer them; I, the God of Israel, will not forsake them.
ISA|41|18|I will make rivers flow on barren heights, and springs within the valleys. I will turn the desert into pools of water, and the parched ground into springs.
ISA|41|19|I will put in the desert the cedar and the acacia, the myrtle and the olive. I will set pines in the wasteland, the fir and the cypress together,
ISA|41|20|so that people may see and know, may consider and understand, that the hand of the LORD has done this, that the Holy One of Israel has created it.
ISA|41|21|"Present your case," says the LORD. "Set forth your arguments," says Jacob's King.
ISA|41|22|"Bring in your idols to tell us what is going to happen. Tell us what the former things were, so that we may consider them and know their final outcome. Or declare to us the things to come,
ISA|41|23|tell us what the future holds, so we may know that you are gods. Do something, whether good or bad, so that we will be dismayed and filled with fear.
ISA|41|24|But you are less than nothing and your works are utterly worthless; he who chooses you is detestable.
ISA|41|25|"I have stirred up one from the north, and he comes- one from the rising sun who calls on my name. He treads on rulers as if they were mortar, as if he were a potter treading the clay.
ISA|41|26|Who told of this from the beginning, so we could know, or beforehand, so we could say, 'He was right'? No one told of this, no one foretold it, no one heard any words from you.
ISA|41|27|I was the first to tell Zion, 'Look, here they are!' I gave to Jerusalem a messenger of good tidings.
ISA|41|28|I look but there is no one- no one among them to give counsel, no one to give answer when I ask them.
ISA|41|29|See, they are all false! Their deeds amount to nothing; their images are but wind and confusion.
ISA|42|1|"Here is my servant, whom I uphold, my chosen one in whom I delight; I will put my Spirit on him and he will bring justice to the nations.
ISA|42|2|He will not shout or cry out, or raise his voice in the streets.
ISA|42|3|A bruised reed he will not break, and a smoldering wick he will not snuff out. In faithfulness he will bring forth justice;
ISA|42|4|he will not falter or be discouraged till he establishes justice on earth. In his law the islands will put their hope."
ISA|42|5|This is what God the LORD says- he who created the heavens and stretched them out, who spread out the earth and all that comes out of it, who gives breath to its people, and life to those who walk on it:
ISA|42|6|"I, the LORD, have called you in righteousness; I will take hold of your hand. I will keep you and will make you to be a covenant for the people and a light for the Gentiles,
ISA|42|7|to open eyes that are blind, to free captives from prison and to release from the dungeon those who sit in darkness.
ISA|42|8|"I am the LORD; that is my name! I will not give my glory to another or my praise to idols.
ISA|42|9|See, the former things have taken place, and new things I declare; before they spring into being I announce them to you."
ISA|42|10|Sing to the LORD a new song, his praise from the ends of the earth, you who go down to the sea, and all that is in it, you islands, and all who live in them.
ISA|42|11|Let the desert and its towns raise their voices; let the settlements where Kedar lives rejoice. Let the people of Sela sing for joy; let them shout from the mountaintops.
ISA|42|12|Let them give glory to the LORD and proclaim his praise in the islands.
ISA|42|13|The LORD will march out like a mighty man, like a warrior he will stir up his zeal; with a shout he will raise the battle cry and will triumph over his enemies.
ISA|42|14|"For a long time I have kept silent, I have been quiet and held myself back. But now, like a woman in childbirth, I cry out, I gasp and pant.
ISA|42|15|I will lay waste the mountains and hills and dry up all their vegetation; I will turn rivers into islands and dry up the pools.
ISA|42|16|I will lead the blind by ways they have not known, along unfamiliar paths I will guide them; I will turn the darkness into light before them and make the rough places smooth. These are the things I will do; I will not forsake them.
ISA|42|17|But those who trust in idols, who say to images, 'You are our gods,' will be turned back in utter shame.
ISA|42|18|"Hear, you deaf; look, you blind, and see!
ISA|42|19|Who is blind but my servant, and deaf like the messenger I send? Who is blind like the one committed to me, blind like the servant of the LORD?
ISA|42|20|You have seen many things, but have paid no attention; your ears are open, but you hear nothing."
ISA|42|21|It pleased the LORD for the sake of his righteousness to make his law great and glorious.
ISA|42|22|But this is a people plundered and looted, all of them trapped in pits or hidden away in prisons. They have become plunder, with no one to rescue them; they have been made loot, with no one to say, "Send them back."
ISA|42|23|Which of you will listen to this or pay close attention in time to come?
ISA|42|24|Who handed Jacob over to become loot, and Israel to the plunderers? Was it not the LORD, against whom we have sinned? For they would not follow his ways; they did not obey his law.
ISA|42|25|So he poured out on them his burning anger, the violence of war. It enveloped them in flames, yet they did not understand; it consumed them, but they did not take it to heart.
ISA|43|1|But now, this is what the LORD says- he who created you, O Jacob, he who formed you, O Israel: "Fear not, for I have redeemed you; I have summoned you by name; you are mine.
ISA|43|2|When you pass through the waters, I will be with you; and when you pass through the rivers, they will not sweep over you. When you walk through the fire, you will not be burned; the flames will not set you ablaze.
ISA|43|3|For I am the LORD, your God, the Holy One of Israel, your Savior; I give Egypt for your ransom, Cush and Seba in your stead.
ISA|43|4|Since you are precious and honored in my sight, and because I love you, I will give men in exchange for you, and people in exchange for your life.
ISA|43|5|Do not be afraid, for I am with you; I will bring your children from the east and gather you from the west.
ISA|43|6|I will say to the north, 'Give them up!' and to the south, 'Do not hold them back.' Bring my sons from afar and my daughters from the ends of the earth-
ISA|43|7|everyone who is called by my name, whom I created for my glory, whom I formed and made."
ISA|43|8|Lead out those who have eyes but are blind, who have ears but are deaf.
ISA|43|9|All the nations gather together and the peoples assemble. Which of them foretold this and proclaimed to us the former things? Let them bring in their witnesses to prove they were right, so that others may hear and say, "It is true."
ISA|43|10|"You are my witnesses," declares the LORD, "and my servant whom I have chosen, so that you may know and believe me and understand that I am he. Before me no god was formed, nor will there be one after me.
ISA|43|11|I, even I, am the LORD, and apart from me there is no savior.
ISA|43|12|I have revealed and saved and proclaimed- I, and not some foreign god among you. You are my witnesses," declares the LORD, "that I am God.
ISA|43|13|Yes, and from ancient days I am he. No one can deliver out of my hand. When I act, who can reverse it?"
ISA|43|14|This is what the LORD says- your Redeemer, the Holy One of Israel: "For your sake I will send to Babylon and bring down as fugitives all the Babylonians, in the ships in which they took pride.
ISA|43|15|I am the LORD, your Holy One, Israel's Creator, your King."
ISA|43|16|This is what the LORD says- he who made a way through the sea, a path through the mighty waters,
ISA|43|17|who drew out the chariots and horses, the army and reinforcements together, and they lay there, never to rise again, extinguished, snuffed out like a wick:
ISA|43|18|"Forget the former things; do not dwell on the past.
ISA|43|19|See, I am doing a new thing! Now it springs up; do you not perceive it? I am making a way in the desert and streams in the wasteland.
ISA|43|20|The wild animals honor me, the jackals and the owls, because I provide water in the desert and streams in the wasteland, to give drink to my people, my chosen,
ISA|43|21|the people I formed for myself that they may proclaim my praise.
ISA|43|22|"Yet you have not called upon me, O Jacob, you have not wearied yourselves for me, O Israel.
ISA|43|23|You have not brought me sheep for burnt offerings, nor honored me with your sacrifices. I have not burdened you with grain offerings nor wearied you with demands for incense.
ISA|43|24|You have not bought any fragrant calamus for me, or lavished on me the fat of your sacrifices. But you have burdened me with your sins and wearied me with your offenses.
ISA|43|25|"I, even I, am he who blots out your transgressions, for my own sake, and remembers your sins no more.
ISA|43|26|Review the past for me, let us argue the matter together; state the case for your innocence.
ISA|43|27|Your first father sinned; your spokesmen rebelled against me.
ISA|43|28|So I will disgrace the dignitaries of your temple, and I will consign Jacob to destruction and Israel to scorn.
ISA|44|1|"But now listen, O Jacob, my servant, Israel, whom I have chosen.
ISA|44|2|This is what the LORD says- he who made you, who formed you in the womb, and who will help you: Do not be afraid, O Jacob, my servant, Jeshurun, whom I have chosen.
ISA|44|3|For I will pour water on the thirsty land, and streams on the dry ground; I will pour out my Spirit on your offspring, and my blessing on your descendants.
ISA|44|4|They will spring up like grass in a meadow, like poplar trees by flowing streams.
ISA|44|5|One will say, 'I belong to the LORD '; another will call himself by the name of Jacob; still another will write on his hand, 'The LORD's,' and will take the name Israel.
ISA|44|6|"This is what the LORD says- Israel's King and Redeemer, the LORD Almighty: I am the first and I am the last; apart from me there is no God.
ISA|44|7|Who then is like me? Let him proclaim it. Let him declare and lay out before me what has happened since I established my ancient people, and what is yet to come- yes, let him foretell what will come.
ISA|44|8|Do not tremble, do not be afraid. Did I not proclaim this and foretell it long ago? You are my witnesses. Is there any God besides me? No, there is no other Rock; I know not one."
ISA|44|9|All who make idols are nothing, and the things they treasure are worthless. Those who would speak up for them are blind; they are ignorant, to their own shame.
ISA|44|10|Who shapes a god and casts an idol, which can profit him nothing?
ISA|44|11|He and his kind will be put to shame; craftsmen are nothing but men. Let them all come together and take their stand; they will be brought down to terror and infamy.
ISA|44|12|The blacksmith takes a tool and works with it in the coals; he shapes an idol with hammers, he forges it with the might of his arm. He gets hungry and loses his strength; he drinks no water and grows faint.
ISA|44|13|The carpenter measures with a line and makes an outline with a marker; he roughs it out with chisels and marks it with compasses. He shapes it in the form of man, of man in all his glory, that it may dwell in a shrine.
ISA|44|14|He cut down cedars, or perhaps took a cypress or oak. He let it grow among the trees of the forest, or planted a pine, and the rain made it grow.
ISA|44|15|It is man's fuel for burning; some of it he takes and warms himself, he kindles a fire and bakes bread. But he also fashions a god and worships it; he makes an idol and bows down to it.
ISA|44|16|Half of the wood he burns in the fire; over it he prepares his meal, he roasts his meat and eats his fill. He also warms himself and says, "Ah! I am warm; I see the fire."
ISA|44|17|From the rest he makes a god, his idol; he bows down to it and worships. He prays to it and says, "Save me; you are my god."
ISA|44|18|They know nothing, they understand nothing; their eyes are plastered over so they cannot see, and their minds closed so they cannot understand.
ISA|44|19|No one stops to think, no one has the knowledge or understanding to say, "Half of it I used for fuel; I even baked bread over its coals, I roasted meat and I ate. Shall I make a detestable thing from what is left? Shall I bow down to a block of wood?"
ISA|44|20|He feeds on ashes, a deluded heart misleads him; he cannot save himself, or say, "Is not this thing in my right hand a lie?"
ISA|44|21|"Remember these things, O Jacob, for you are my servant, O Israel. I have made you, you are my servant; O Israel, I will not forget you.
ISA|44|22|I have swept away your offenses like a cloud, your sins like the morning mist. Return to me, for I have redeemed you."
ISA|44|23|Sing for joy, O heavens, for the LORD has done this; shout aloud, O earth beneath. Burst into song, you mountains, you forests and all your trees, for the LORD has redeemed Jacob, he displays his glory in Israel.
ISA|44|24|"This is what the LORD says- your Redeemer, who formed you in the womb: I am the LORD, who has made all things, who alone stretched out the heavens, who spread out the earth by myself,
ISA|44|25|who foils the signs of false prophets and makes fools of diviners, who overthrows the learning of the wise and turns it into nonsense,
ISA|44|26|who carries out the words of his servants and fulfills the predictions of his messengers, who says of Jerusalem, 'It shall be inhabited,' of the towns of Judah, 'They shall be built,' and of their ruins, 'I will restore them,'
ISA|44|27|who says to the watery deep, 'Be dry, and I will dry up your streams,'
ISA|44|28|who says of Cyrus, 'He is my shepherd and will accomplish all that I please; he will say of Jerusalem, "Let it be rebuilt," and of the temple, "Let its foundations be laid."'
ISA|45|1|"This is what the LORD says to his anointed, to Cyrus, whose right hand I take hold of to subdue nations before him and to strip kings of their armor, to open doors before him so that gates will not be shut:
ISA|45|2|I will go before you and will level the mountains; I will break down gates of bronze and cut through bars of iron.
ISA|45|3|I will give you the treasures of darkness, riches stored in secret places, so that you may know that I am the LORD, the God of Israel, who summons you by name.
ISA|45|4|For the sake of Jacob my servant, of Israel my chosen, I summon you by name and bestow on you a title of honor, though you do not acknowledge me.
ISA|45|5|I am the LORD, and there is no other; apart from me there is no God. I will strengthen you, though you have not acknowledged me,
ISA|45|6|so that from the rising of the sun to the place of its setting men may know there is none besides me. I am the LORD, and there is no other.
ISA|45|7|I form the light and create darkness, I bring prosperity and create disaster; I, the LORD, do all these things.
ISA|45|8|"You heavens above, rain down righteousness; let the clouds shower it down. Let the earth open wide, let salvation spring up, let righteousness grow with it; I, the LORD, have created it.
ISA|45|9|"Woe to him who quarrels with his Maker, to him who is but a potsherd among the potsherds on the ground. Does the clay say to the potter, 'What are you making?' Does your work say, 'He has no hands'?
ISA|45|10|Woe to him who says to his father, 'What have you begotten?' or to his mother, 'What have you brought to birth?'
ISA|45|11|"This is what the LORD says- the Holy One of Israel, and its Maker: Concerning things to come, do you question me about my children, or give me orders about the work of my hands?
ISA|45|12|It is I who made the earth and created mankind upon it. My own hands stretched out the heavens; I marshaled their starry hosts.
ISA|45|13|I will raise up Cyrus in my righteousness: I will make all his ways straight. He will rebuild my city and set my exiles free, but not for a price or reward, says the LORD Almighty."
ISA|45|14|This is what the LORD says: "The products of Egypt and the merchandise of Cush, and those tall Sabeans- they will come over to you and will be yours; they will trudge behind you, coming over to you in chains. They will bow down before you and plead with you, saying, 'Surely God is with you, and there is no other; there is no other god.'"
ISA|45|15|Truly you are a God who hides himself, O God and Savior of Israel.
ISA|45|16|All the makers of idols will be put to shame and disgraced; they will go off into disgrace together.
ISA|45|17|But Israel will be saved by the LORD with an everlasting salvation; you will never be put to shame or disgraced, to ages everlasting.
ISA|45|18|For this is what the LORD says- he who created the heavens, he is God; he who fashioned and made the earth, he founded it; he did not create it to be empty, but formed it to be inhabited- he says: "I am the LORD, and there is no other.
ISA|45|19|I have not spoken in secret, from somewhere in a land of darkness; I have not said to Jacob's descendants, 'Seek me in vain.' I, the LORD, speak the truth; I declare what is right.
ISA|45|20|"Gather together and come; assemble, you fugitives from the nations. Ignorant are those who carry about idols of wood, who pray to gods that cannot save.
ISA|45|21|Declare what is to be, present it- let them take counsel together. Who foretold this long ago, who declared it from the distant past? Was it not I, the LORD? And there is no God apart from me, a righteous God and a Savior; there is none but me.
ISA|45|22|"Turn to me and be saved, all you ends of the earth; for I am God, and there is no other.
ISA|45|23|By myself I have sworn, my mouth has uttered in all integrity a word that will not be revoked: Before me every knee will bow; by me every tongue will swear.
ISA|45|24|They will say of me, 'In the LORD alone are righteousness and strength.'" All who have raged against him will come to him and be put to shame.
ISA|45|25|But in the LORD all the descendants of Israel will be found righteous and will exult.
ISA|46|1|Bel bows down, Nebo stoops low; their idols are borne by beasts of burden. The images that are carried about are burdensome, a burden for the weary.
ISA|46|2|They stoop and bow down together; unable to rescue the burden, they themselves go off into captivity.
ISA|46|3|"Listen to me, O house of Jacob, all you who remain of the house of Israel, you whom I have upheld since you were conceived, and have carried since your birth.
ISA|46|4|Even to your old age and gray hairs I am he, I am he who will sustain you. I have made you and I will carry you; I will sustain you and I will rescue you.
ISA|46|5|"To whom will you compare me or count me equal? To whom will you liken me that we may be compared?
ISA|46|6|Some pour out gold from their bags and weigh out silver on the scales; they hire a goldsmith to make it into a god, and they bow down and worship it.
ISA|46|7|They lift it to their shoulders and carry it; they set it up in its place, and there it stands. From that spot it cannot move. Though one cries out to it, it does not answer; it cannot save him from his troubles.
ISA|46|8|"Remember this, fix it in mind, take it to heart, you rebels.
ISA|46|9|Remember the former things, those of long ago; I am God, and there is no other; I am God, and there is none like me.
ISA|46|10|I make known the end from the beginning, from ancient times, what is still to come. I say: My purpose will stand, and I will do all that I please.
ISA|46|11|From the east I summon a bird of prey; from a far-off land, a man to fulfill my purpose. What I have said, that will I bring about; what I have planned, that will I do.
ISA|46|12|Listen to me, you stubborn-hearted, you who are far from righteousness.
ISA|46|13|I am bringing my righteousness near, it is not far away; and my salvation will not be delayed. I will grant salvation to Zion, my splendor to Israel.
ISA|47|1|"Go down, sit in the dust, Virgin Daughter of Babylon; sit on the ground without a throne, Daughter of the Babylonians. No more will you be called tender or delicate.
ISA|47|2|Take millstones and grind flour; take off your veil. Lift up your skirts, bare your legs, and wade through the streams.
ISA|47|3|Your nakedness will be exposed and your shame uncovered. I will take vengeance; I will spare no one."
ISA|47|4|Our Redeemer-the LORD Almighty is his name- is the Holy One of Israel.
ISA|47|5|"Sit in silence, go into darkness, Daughter of the Babylonians; no more will you be called queen of kingdoms.
ISA|47|6|I was angry with my people and desecrated my inheritance; I gave them into your hand, and you showed them no mercy. Even on the aged you laid a very heavy yoke.
ISA|47|7|You said, 'I will continue forever- the eternal queen!' But you did not consider these things or reflect on what might happen.
ISA|47|8|"Now then, listen, you wanton creature, lounging in your security and saying to yourself, 'I am, and there is none besides me. I will never be a widow or suffer the loss of children.'
ISA|47|9|Both of these will overtake you in a moment, on a single day: loss of children and widowhood. They will come upon you in full measure, in spite of your many sorceries and all your potent spells.
ISA|47|10|You have trusted in your wickedness and have said, 'No one sees me.' Your wisdom and knowledge mislead you when you say to yourself, 'I am, and there is none besides me.'
ISA|47|11|Disaster will come upon you, and you will not know how to conjure it away. A calamity will fall upon you that you cannot ward off with a ransom; a catastrophe you cannot foresee will suddenly come upon you.
ISA|47|12|"Keep on, then, with your magic spells and with your many sorceries, which you have labored at since childhood. Perhaps you will succeed, perhaps you will cause terror.
ISA|47|13|All the counsel you have received has only worn you out! Let your astrologers come forward, those stargazers who make predictions month by month, let them save you from what is coming upon you.
ISA|47|14|Surely they are like stubble; the fire will burn them up. They cannot even save themselves from the power of the flame. Here are no coals to warm anyone; here is no fire to sit by.
ISA|47|15|That is all they can do for you- these you have labored with and trafficked with since childhood. Each of them goes on in his error; there is not one that can save you.
ISA|48|1|"Listen to this, O house of Jacob, you who are called by the name of Israel and come from the line of Judah, you who take oaths in the name of the LORD and invoke the God of Israel- but not in truth or righteousness-
ISA|48|2|you who call yourselves citizens of the holy city and rely on the God of Israel- the LORD Almighty is his name:
ISA|48|3|I foretold the former things long ago, my mouth announced them and I made them known; then suddenly I acted, and they came to pass.
ISA|48|4|For I knew how stubborn you were; the sinews of your neck were iron, your forehead was bronze.
ISA|48|5|Therefore I told you these things long ago; before they happened I announced them to you so that you could not say, 'My idols did them; my wooden image and metal god ordained them.'
ISA|48|6|You have heard these things; look at them all. Will you not admit them? "From now on I will tell you of new things, of hidden things unknown to you.
ISA|48|7|They are created now, and not long ago; you have not heard of them before today. So you cannot say, 'Yes, I knew of them.'
ISA|48|8|You have neither heard nor understood; from of old your ear has not been open. Well do I know how treacherous you are; you were called a rebel from birth.
ISA|48|9|For my own name's sake I delay my wrath; for the sake of my praise I hold it back from you, so as not to cut you off.
ISA|48|10|See, I have refined you, though not as silver; I have tested you in the furnace of affliction.
ISA|48|11|For my own sake, for my own sake, I do this. How can I let myself be defamed? I will not yield my glory to another.
ISA|48|12|"Listen to me, O Jacob, Israel, whom I have called: I am he; I am the first and I am the last.
ISA|48|13|My own hand laid the foundations of the earth, and my right hand spread out the heavens; when I summon them, they all stand up together.
ISA|48|14|"Come together, all of you, and listen: Which of the idols has foretold these things? The LORD's chosen ally will carry out his purpose against Babylon; his arm will be against the Babylonians.
ISA|48|15|I, even I, have spoken; yes, I have called him. I will bring him, and he will succeed in his mission.
ISA|48|16|"Come near me and listen to this: "From the first announcement I have not spoken in secret; at the time it happens, I am there." And now the Sovereign LORD has sent me, with his Spirit.
ISA|48|17|This is what the LORD says- your Redeemer, the Holy One of Israel: "I am the LORD your God, who teaches you what is best for you, who directs you in the way you should go.
ISA|48|18|If only you had paid attention to my commands, your peace would have been like a river, your righteousness like the waves of the sea.
ISA|48|19|Your descendants would have been like the sand, your children like its numberless grains; their name would never be cut off nor destroyed from before me."
ISA|48|20|Leave Babylon, flee from the Babylonians! Announce this with shouts of joy and proclaim it. Send it out to the ends of the earth; say, "The LORD has redeemed his servant Jacob."
ISA|48|21|They did not thirst when he led them through the deserts; he made water flow for them from the rock; he split the rock and water gushed out.
ISA|48|22|"There is no peace," says the LORD, "for the wicked."
ISA|49|1|Listen to me, you islands; hear this, you distant nations: Before I was born the LORD called me; from my birth he has made mention of my name.
ISA|49|2|He made my mouth like a sharpened sword, in the shadow of his hand he hid me; he made me into a polished arrow and concealed me in his quiver.
ISA|49|3|He said to me, "You are my servant, Israel, in whom I will display my splendor."
ISA|49|4|But I said, "I have labored to no purpose; I have spent my strength in vain and for nothing. Yet what is due me is in the LORD's hand, and my reward is with my God."
ISA|49|5|And now the LORD says- he who formed me in the womb to be his servant to bring Jacob back to him and gather Israel to himself, for I am honored in the eyes of the LORD and my God has been my strength-
ISA|49|6|he says: "It is too small a thing for you to be my servant to restore the tribes of Jacob and bring back those of Israel I have kept. I will also make you a light for the Gentiles, that you may bring my salvation to the ends of the earth."
ISA|49|7|This is what the LORD says- the Redeemer and Holy One of Israel- to him who was despised and abhorred by the nation, to the servant of rulers: "Kings will see you and rise up, princes will see and bow down, because of the LORD, who is faithful, the Holy One of Israel, who has chosen you."
ISA|49|8|This is what the LORD says: "In the time of my favor I will answer you, and in the day of salvation I will help you; I will keep you and will make you to be a covenant for the people, to restore the land and to reassign its desolate inheritances,
ISA|49|9|to say to the captives, 'Come out,' and to those in darkness, 'Be free!'"They will feed beside the roads and find pasture on every barren hill.
ISA|49|10|They will neither hunger nor thirst, nor will the desert heat or the sun beat upon them. He who has compassion on them will guide them and lead them beside springs of water.
ISA|49|11|I will turn all my mountains into roads, and my highways will be raised up.
ISA|49|12|See, they will come from afar- some from the north, some from the west, some from the region of Aswan. "
ISA|49|13|Shout for joy, O heavens; rejoice, O earth; burst into song, O mountains! For the LORD comforts his people and will have compassion on his afflicted ones.
ISA|49|14|But Zion said, "The LORD has forsaken me, the Lord has forgotten me."
ISA|49|15|"Can a mother forget the baby at her breast and have no compassion on the child she has borne? Though she may forget, I will not forget you!
ISA|49|16|See, I have engraved you on the palms of my hands; your walls are ever before me.
ISA|49|17|Your sons hasten back, and those who laid you waste depart from you.
ISA|49|18|Lift up your eyes and look around; all your sons gather and come to you. As surely as I live," declares the LORD, "you will wear them all as ornaments; you will put them on, like a bride.
ISA|49|19|"Though you were ruined and made desolate and your land laid waste, now you will be too small for your people, and those who devoured you will be far away.
ISA|49|20|The children born during your bereavement will yet say in your hearing, 'This place is too small for us; give us more space to live in.'
ISA|49|21|Then you will say in your heart, 'Who bore me these? I was bereaved and barren; I was exiled and rejected. Who brought these up? I was left all alone, but these-where have they come from?'"
ISA|49|22|This is what the Sovereign LORD says: "See, I will beckon to the Gentiles, I will lift up my banner to the peoples; they will bring your sons in their arms and carry your daughters on their shoulders.
ISA|49|23|Kings will be your foster fathers, and their queens your nursing mothers. They will bow down before you with their faces to the ground; they will lick the dust at your feet. Then you will know that I am the LORD; those who hope in me will not be disappointed."
ISA|49|24|Can plunder be taken from warriors, or captives rescued from the fierce?
ISA|49|25|But this is what the LORD says: "Yes, captives will be taken from warriors, and plunder retrieved from the fierce; I will contend with those who contend with you, and your children I will save.
ISA|49|26|I will make your oppressors eat their own flesh; they will be drunk on their own blood, as with wine. Then all mankind will know that I, the LORD, am your Savior, your Redeemer, the Mighty One of Jacob."
ISA|50|1|This is what the LORD says: "Where is your mother's certificate of divorce with which I sent her away? Or to which of my creditors did I sell you? Because of your sins you were sold; because of your transgressions your mother was sent away.
ISA|50|2|When I came, why was there no one? When I called, why was there no one to answer? Was my arm too short to ransom you? Do I lack the strength to rescue you? By a mere rebuke I dry up the sea, I turn rivers into a desert; their fish rot for lack of water and die of thirst.
ISA|50|3|I clothe the sky with darkness and make sackcloth its covering."
ISA|50|4|The Sovereign LORD has given me an instructed tongue, to know the word that sustains the weary. He wakens me morning by morning, wakens my ear to listen like one being taught.
ISA|50|5|The Sovereign LORD has opened my ears, and I have not been rebellious; I have not drawn back.
ISA|50|6|I offered my back to those who beat me, my cheeks to those who pulled out my beard; I did not hide my face from mocking and spitting.
ISA|50|7|Because the Sovereign LORD helps me, I will not be disgraced. Therefore have I set my face like flint, and I know I will not be put to shame.
ISA|50|8|He who vindicates me is near. Who then will bring charges against me? Let us face each other! Who is my accuser? Let him confront me!
ISA|50|9|It is the Sovereign LORD who helps me. Who is he that will condemn me? They will all wear out like a garment; the moths will eat them up.
ISA|50|10|Who among you fears the LORD and obeys the word of his servant? Let him who walks in the dark, who has no light, trust in the name of the LORD and rely on his God.
ISA|50|11|But now, all you who light fires and provide yourselves with flaming torches, go, walk in the light of your fires and of the torches you have set ablaze. This is what you shall receive from my hand: You will lie down in torment.
ISA|51|1|"Listen to me, you who pursue righteousness and who seek the LORD: Look to the rock from which you were cut and to the quarry from which you were hewn;
ISA|51|2|look to Abraham, your father, and to Sarah, who gave you birth. When I called him he was but one, and I blessed him and made him many.
ISA|51|3|The LORD will surely comfort Zion and will look with compassion on all her ruins; he will make her deserts like Eden, her wastelands like the garden of the LORD. Joy and gladness will be found in her, thanksgiving and the sound of singing.
ISA|51|4|"Listen to me, my people; hear me, my nation: The law will go out from me; my justice will become a light to the nations.
ISA|51|5|My righteousness draws near speedily, my salvation is on the way, and my arm will bring justice to the nations. The islands will look to me and wait in hope for my arm.
ISA|51|6|Lift up your eyes to the heavens, look at the earth beneath; the heavens will vanish like smoke, the earth will wear out like a garment and its inhabitants die like flies. But my salvation will last forever, my righteousness will never fail.
ISA|51|7|"Hear me, you who know what is right, you people who have my law in your hearts: Do not fear the reproach of men or be terrified by their insults.
ISA|51|8|For the moth will eat them up like a garment; the worm will devour them like wool. But my righteousness will last forever, my salvation through all generations."
ISA|51|9|Awake, awake! Clothe yourself with strength, O arm of the LORD; awake, as in days gone by, as in generations of old. Was it not you who cut Rahab to pieces, who pierced that monster through?
ISA|51|10|Was it not you who dried up the sea, the waters of the great deep, who made a road in the depths of the sea so that the redeemed might cross over?
ISA|51|11|The ransomed of the LORD will return. They will enter Zion with singing; everlasting joy will crown their heads. Gladness and joy will overtake them, and sorrow and sighing will flee away.
ISA|51|12|"I, even I, am he who comforts you. Who are you that you fear mortal men, the sons of men, who are but grass,
ISA|51|13|that you forget the LORD your Maker, who stretched out the heavens and laid the foundations of the earth, that you live in constant terror every day because of the wrath of the oppressor, who is bent on destruction? For where is the wrath of the oppressor?
ISA|51|14|The cowering prisoners will soon be set free; they will not die in their dungeon, nor will they lack bread.
ISA|51|15|For I am the LORD your God, who churns up the sea so that its waves roar- the LORD Almighty is his name.
ISA|51|16|I have put my words in your mouth and covered you with the shadow of my hand- I who set the heavens in place, who laid the foundations of the earth, and who say to Zion, 'You are my people.'"
ISA|51|17|Awake, awake! Rise up, O Jerusalem, you who have drunk from the hand of the LORD the cup of his wrath, you who have drained to its dregs the goblet that makes men stagger.
ISA|51|18|Of all the sons she bore there was none to guide her; of all the sons she reared there was none to take her by the hand.
ISA|51|19|These double calamities have come upon you- who can comfort you?- ruin and destruction, famine and sword- who can console you?
ISA|51|20|Your sons have fainted; they lie at the head of every street, like antelope caught in a net. They are filled with the wrath of the LORD and the rebuke of your God.
ISA|51|21|Therefore hear this, you afflicted one, made drunk, but not with wine.
ISA|51|22|This is what your Sovereign LORD says, your God, who defends his people: "See, I have taken out of your hand the cup that made you stagger; from that cup, the goblet of my wrath, you will never drink again.
ISA|51|23|I will put it into the hands of your tormentors, who said to you, 'Fall prostrate that we may walk over you.' And you made your back like the ground, like a street to be walked over."
ISA|52|1|Awake, awake, O Zion, clothe yourself with strength. Put on your garments of splendor, O Jerusalem, the holy city. The uncircumcised and defiled will not enter you again.
ISA|52|2|Shake off your dust; rise up, sit enthroned, O Jerusalem. Free yourself from the chains on your neck, O captive Daughter of Zion.
ISA|52|3|For this is what the LORD says: "You were sold for nothing, and without money you will be redeemed."
ISA|52|4|For this is what the Sovereign LORD says: "At first my people went down to Egypt to live; lately, Assyria has oppressed them.
ISA|52|5|"And now what do I have here?" declares the LORD. "For my people have been taken away for nothing, and those who rule them mock, "declares the LORD. "And all day long my name is constantly blasphemed.
ISA|52|6|Therefore my people will know my name; therefore in that day they will know that it is I who foretold it. Yes, it is I."
ISA|52|7|How beautiful on the mountains are the feet of those who bring good news, who proclaim peace, who bring good tidings, who proclaim salvation, who say to Zion, "Your God reigns!"
ISA|52|8|Listen! Your watchmen lift up their voices; together they shout for joy. When the LORD returns to Zion, they will see it with their own eyes.
ISA|52|9|Burst into songs of joy together, you ruins of Jerusalem, for the LORD has comforted his people, he has redeemed Jerusalem.
ISA|52|10|The LORD will lay bare his holy arm in the sight of all the nations, and all the ends of the earth will see the salvation of our God.
ISA|52|11|Depart, depart, go out from there! Touch no unclean thing! Come out from it and be pure, you who carry the vessels of the LORD.
ISA|52|12|But you will not leave in haste or go in flight; for the LORD will go before you, the God of Israel will be your rear guard.
ISA|52|13|See, my servant will act wisely; he will be raised and lifted up and highly exalted.
ISA|52|14|Just as there were many who were appalled at him - his appearance was so disfigured beyond that of any man and his form marred beyond human likeness-
ISA|52|15|so will he sprinkle many nations, and kings will shut their mouths because of him. For what they were not told, they will see, and what they have not heard, they will understand.
ISA|53|1|Who has believed our message and to whom has the arm of the LORD been revealed?
ISA|53|2|He grew up before him like a tender shoot, and like a root out of dry ground. He had no beauty or majesty to attract us to him, nothing in his appearance that we should desire him.
ISA|53|3|He was despised and rejected by men, a man of sorrows, and familiar with suffering. Like one from whom men hide their faces he was despised, and we esteemed him not.
ISA|53|4|Surely he took up our infirmities and carried our sorrows, yet we considered him stricken by God, smitten by him, and afflicted.
ISA|53|5|But he was pierced for our transgressions, he was crushed for our iniquities; the punishment that brought us peace was upon him, and by his wounds we are healed.
ISA|53|6|We all, like sheep, have gone astray, each of us has turned to his own way; and the LORD has laid on him the iniquity of us all.
ISA|53|7|He was oppressed and afflicted, yet he did not open his mouth; he was led like a lamb to the slaughter, and as a sheep before her shearers is silent, so he did not open his mouth.
ISA|53|8|By oppression and judgment he was taken away. And who can speak of his descendants? For he was cut off from the land of the living; for the transgression of my people he was stricken.
ISA|53|9|He was assigned a grave with the wicked, and with the rich in his death, though he had done no violence, nor was any deceit in his mouth.
ISA|53|10|Yet it was the LORD's will to crush him and cause him to suffer, and though the LORD makes his life a guilt offering, he will see his offspring and prolong his days, and the will of the LORD will prosper in his hand.
ISA|53|11|After the suffering of his soul, he will see the light of life and be satisfied; by his knowledge my righteous servant will justify many, and he will bear their iniquities.
ISA|53|12|Therefore I will give him a portion among the great, and he will divide the spoils with the strong, because he poured out his life unto death, and was numbered with the transgressors. For he bore the sin of many, and made intercession for the transgressors.
ISA|54|1|"Sing, O barren woman, you who never bore a child; burst into song, shout for joy, you who were never in labor; because more are the children of the desolate woman than of her who has a husband," says the LORD.
ISA|54|2|"Enlarge the place of your tent, stretch your tent curtains wide, do not hold back; lengthen your cords, strengthen your stakes.
ISA|54|3|For you will spread out to the right and to the left; your descendants will dispossess nations and settle in their desolate cities.
ISA|54|4|"Do not be afraid; you will not suffer shame. Do not fear disgrace; you will not be humiliated. You will forget the shame of your youth and remember no more the reproach of your widowhood.
ISA|54|5|For your Maker is your husband- the LORD Almighty is his name- the Holy One of Israel is your Redeemer; he is called the God of all the earth.
ISA|54|6|The LORD will call you back as if you were a wife deserted and distressed in spirit- a wife who married young, only to be rejected," says your God.
ISA|54|7|"For a brief moment I abandoned you, but with deep compassion I will bring you back.
ISA|54|8|In a surge of anger I hid my face from you for a moment, but with everlasting kindness I will have compassion on you," says the LORD your Redeemer.
ISA|54|9|"To me this is like the days of Noah, when I swore that the waters of Noah would never again cover the earth. So now I have sworn not to be angry with you, never to rebuke you again.
ISA|54|10|Though the mountains be shaken and the hills be removed, yet my unfailing love for you will not be shaken nor my covenant of peace be removed," says the LORD, who has compassion on you.
ISA|54|11|"O afflicted city, lashed by storms and not comforted, I will build you with stones of turquoise, your foundations with sapphires.
ISA|54|12|I will make your battlements of rubies, your gates of sparkling jewels, and all your walls of precious stones.
ISA|54|13|All your sons will be taught by the LORD, and great will be your children's peace.
ISA|54|14|In righteousness you will be established: Tyranny will be far from you; you will have nothing to fear. Terror will be far removed; it will not come near you.
ISA|54|15|If anyone does attack you, it will not be my doing; whoever attacks you will surrender to you.
ISA|54|16|"See, it is I who created the blacksmith who fans the coals into flame and forges a weapon fit for its work. And it is I who have created the destroyer to work havoc;
ISA|54|17|no weapon forged against you will prevail, and you will refute every tongue that accuses you. This is the heritage of the servants of the LORD, and this is their vindication from me," declares the LORD.
ISA|55|1|"Come, all you who are thirsty, come to the waters; and you who have no money, come, buy and eat! Come, buy wine and milk without money and without cost.
ISA|55|2|Why spend money on what is not bread, and your labor on what does not satisfy? Listen, listen to me, and eat what is good, and your soul will delight in the richest of fare.
ISA|55|3|Give ear and come to me; hear me, that your soul may live. I will make an everlasting covenant with you, my faithful love promised to David.
ISA|55|4|See, I have made him a witness to the peoples, a leader and commander of the peoples.
ISA|55|5|Surely you will summon nations you know not, and nations that do not know you will hasten to you, because of the LORD your God, the Holy One of Israel, for he has endowed you with splendor."
ISA|55|6|Seek the LORD while he may be found; call on him while he is near.
ISA|55|7|Let the wicked forsake his way and the evil man his thoughts. Let him turn to the LORD, and he will have mercy on him, and to our God, for he will freely pardon.
ISA|55|8|"For my thoughts are not your thoughts, neither are your ways my ways," declares the LORD.
ISA|55|9|"As the heavens are higher than the earth, so are my ways higher than your ways and my thoughts than your thoughts.
ISA|55|10|As the rain and the snow come down from heaven, and do not return to it without watering the earth and making it bud and flourish, so that it yields seed for the sower and bread for the eater,
ISA|55|11|so is my word that goes out from my mouth: It will not return to me empty, but will accomplish what I desire and achieve the purpose for which I sent it.
ISA|55|12|You will go out in joy and be led forth in peace; the mountains and hills will burst into song before you, and all the trees of the field will clap their hands.
ISA|55|13|Instead of the thornbush will grow the pine tree, and instead of briers the myrtle will grow. This will be for the LORD's renown, for an everlasting sign, which will not be destroyed."
ISA|56|1|This is what the LORD says: "Maintain justice and do what is right, for my salvation is close at hand and my righteousness will soon be revealed.
ISA|56|2|Blessed is the man who does this, the man who holds it fast, who keeps the Sabbath without desecrating it, and keeps his hand from doing any evil."
ISA|56|3|Let no foreigner who has bound himself to the LORD say, "The LORD will surely exclude me from his people." And let not any eunuch complain, "I am only a dry tree."
ISA|56|4|For this is what the LORD says: "To the eunuchs who keep my Sabbaths, who choose what pleases me and hold fast to my covenant-
ISA|56|5|to them I will give within my temple and its walls a memorial and a name better than sons and daughters; I will give them an everlasting name that will not be cut off.
ISA|56|6|And foreigners who bind themselves to the LORD to serve him, to love the name of the LORD, and to worship him, all who keep the Sabbath without desecrating it and who hold fast to my covenant-
ISA|56|7|these I will bring to my holy mountain and give them joy in my house of prayer. Their burnt offerings and sacrifices will be accepted on my altar; for my house will be called a house of prayer for all nations."
ISA|56|8|The Sovereign LORD declares- he who gathers the exiles of Israel: "I will gather still others to them besides those already gathered."
ISA|56|9|Come, all you beasts of the field, come and devour, all you beasts of the forest!
ISA|56|10|Israel's watchmen are blind, they all lack knowledge; they are all mute dogs, they cannot bark; they lie around and dream, they love to sleep.
ISA|56|11|They are dogs with mighty appetites; they never have enough. They are shepherds who lack understanding; they all turn to their own way, each seeks his own gain.
ISA|56|12|"Come," each one cries, "let me get wine! Let us drink our fill of beer! And tomorrow will be like today, or even far better."
ISA|57|1|The righteous perish, and no one ponders it in his heart; devout men are taken away, and no one understands that the righteous are taken away to be spared from evil.
ISA|57|2|Those who walk uprightly enter into peace; they find rest as they lie in death.
ISA|57|3|"But you-come here, you sons of a sorceress, you offspring of adulterers and prostitutes!
ISA|57|4|Whom are you mocking? At whom do you sneer and stick out your tongue? Are you not a brood of rebels, the offspring of liars?
ISA|57|5|You burn with lust among the oaks and under every spreading tree; you sacrifice your children in the ravines and under the overhanging crags.
ISA|57|6|The idols among the smooth stones of the ravines are your portion; they, they are your lot. Yes, to them you have poured out drink offerings and offered grain offerings. In the light of these things, should I relent?
ISA|57|7|You have made your bed on a high and lofty hill; there you went up to offer your sacrifices.
ISA|57|8|Behind your doors and your doorposts you have put your pagan symbols. Forsaking me, you uncovered your bed, you climbed into it and opened it wide; you made a pact with those whose beds you love, and you looked on their nakedness.
ISA|57|9|You went to Molech with olive oil and increased your perfumes. You sent your ambassadors far away; you descended to the grave itself!
ISA|57|10|You were wearied by all your ways, but you would not say, 'It is hopeless.' You found renewal of your strength, and so you did not faint.
ISA|57|11|"Whom have you so dreaded and feared that you have been false to me, and have neither remembered me nor pondered this in your hearts? Is it not because I have long been silent that you do not fear me?
ISA|57|12|I will expose your righteousness and your works, and they will not benefit you.
ISA|57|13|When you cry out for help, let your collection of idols save you! The wind will carry all of them off, a mere breath will blow them away. But the man who makes me his refuge will inherit the land and possess my holy mountain."
ISA|57|14|And it will be said: "Build up, build up, prepare the road! Remove the obstacles out of the way of my people."
ISA|57|15|For this is what the high and lofty One says- he who lives forever, whose name is holy: "I live in a high and holy place, but also with him who is contrite and lowly in spirit, to revive the spirit of the lowly and to revive the heart of the contrite.
ISA|57|16|I will not accuse forever, nor will I always be angry, for then the spirit of man would grow faint before me- the breath of man that I have created.
ISA|57|17|I was enraged by his sinful greed; I punished him, and hid my face in anger, yet he kept on in his willful ways.
ISA|57|18|I have seen his ways, but I will heal him; I will guide him and restore comfort to him,
ISA|57|19|creating praise on the lips of the mourners in Israel. Peace, peace, to those far and near," says the LORD. "And I will heal them."
ISA|57|20|But the wicked are like the tossing sea, which cannot rest, whose waves cast up mire and mud.
ISA|57|21|"There is no peace," says my God, "for the wicked."
ISA|58|1|"Shout it aloud, do not hold back. Raise your voice like a trumpet. Declare to my people their rebellion and to the house of Jacob their sins.
ISA|58|2|For day after day they seek me out; they seem eager to know my ways, as if they were a nation that does what is right and has not forsaken the commands of its God. They ask me for just decisions and seem eager for God to come near them.
ISA|58|3|'Why have we fasted,' they say, 'and you have not seen it? Why have we humbled ourselves, and you have not noticed?'"Yet on the day of your fasting, you do as you please and exploit all your workers.
ISA|58|4|Your fasting ends in quarreling and strife, and in striking each other with wicked fists. You cannot fast as you do today and expect your voice to be heard on high.
ISA|58|5|Is this the kind of fast I have chosen, only a day for a man to humble himself? Is it only for bowing one's head like a reed and for lying on sackcloth and ashes? Is that what you call a fast, a day acceptable to the LORD?
ISA|58|6|"Is not this the kind of fasting I have chosen: to loose the chains of injustice and untie the cords of the yoke, to set the oppressed free and break every yoke?
ISA|58|7|Is it not to share your food with the hungry and to provide the poor wanderer with shelter- when you see the naked, to clothe him, and not to turn away from your own flesh and blood?
ISA|58|8|Then your light will break forth like the dawn, and your healing will quickly appear; then your righteousness will go before you, and the glory of the LORD will be your rear guard.
ISA|58|9|Then you will call, and the LORD will answer; you will cry for help, and he will say: Here am I. "If you do away with the yoke of oppression, with the pointing finger and malicious talk,
ISA|58|10|and if you spend yourselves in behalf of the hungry and satisfy the needs of the oppressed, then your light will rise in the darkness, and your night will become like the noonday.
ISA|58|11|The LORD will guide you always; he will satisfy your needs in a sun-scorched land and will strengthen your frame. You will be like a well-watered garden, like a spring whose waters never fail.
ISA|58|12|Your people will rebuild the ancient ruins and will raise up the age-old foundations; you will be called Repairer of Broken Walls, Restorer of Streets with Dwellings.
ISA|58|13|"If you keep your feet from breaking the Sabbath and from doing as you please on my holy day, if you call the Sabbath a delight and the LORD's holy day honorable, and if you honor it by not going your own way and not doing as you please or speaking idle words,
ISA|58|14|then you will find your joy in the LORD, and I will cause you to ride on the heights of the land and to feast on the inheritance of your father Jacob." The mouth of the LORD has spoken.
ISA|59|1|Surely the arm of the LORD is not too short to save, nor his ear too dull to hear.
ISA|59|2|But your iniquities have separated you from your God; your sins have hidden his face from you, so that he will not hear.
ISA|59|3|For your hands are stained with blood, your fingers with guilt. Your lips have spoken lies, and your tongue mutters wicked things.
ISA|59|4|No one calls for justice; no one pleads his case with integrity. They rely on empty arguments and speak lies; they conceive trouble and give birth to evil.
ISA|59|5|They hatch the eggs of vipers and spin a spider's web. Whoever eats their eggs will die, and when one is broken, an adder is hatched.
ISA|59|6|Their cobwebs are useless for clothing; they cannot cover themselves with what they make. Their deeds are evil deeds, and acts of violence are in their hands.
ISA|59|7|Their feet rush into sin; they are swift to shed innocent blood. Their thoughts are evil thoughts; ruin and destruction mark their ways.
ISA|59|8|The way of peace they do not know; there is no justice in their paths. They have turned them into crooked roads; no one who walks in them will know peace.
ISA|59|9|So justice is far from us, and righteousness does not reach us. We look for light, but all is darkness; for brightness, but we walk in deep shadows.
ISA|59|10|Like the blind we grope along the wall, feeling our way like men without eyes. At midday we stumble as if it were twilight; among the strong, we are like the dead.
ISA|59|11|We all growl like bears; we moan mournfully like doves. We look for justice, but find none; for deliverance, but it is far away.
ISA|59|12|For our offenses are many in your sight, and our sins testify against us. Our offenses are ever with us, and we acknowledge our iniquities:
ISA|59|13|rebellion and treachery against the LORD, turning our backs on our God, fomenting oppression and revolt, uttering lies our hearts have conceived.
ISA|59|14|So justice is driven back, and righteousness stands at a distance; truth has stumbled in the streets, honesty cannot enter.
ISA|59|15|Truth is nowhere to be found, and whoever shuns evil becomes a prey. The LORD looked and was displeased that there was no justice.
ISA|59|16|He saw that there was no one, he was appalled that there was no one to intervene; so his own arm worked salvation for him, and his own righteousness sustained him.
ISA|59|17|He put on righteousness as his breastplate, and the helmet of salvation on his head; he put on the garments of vengeance and wrapped himself in zeal as in a cloak.
ISA|59|18|According to what they have done, so will he repay wrath to his enemies and retribution to his foes; he will repay the islands their due.
ISA|59|19|From the west, men will fear the name of the LORD, and from the rising of the sun, they will revere his glory. For he will come like a pent-up flood that the breath of the LORD drives along.
ISA|59|20|"The Redeemer will come to Zion, to those in Jacob who repent of their sins," declares the LORD.
ISA|59|21|"As for me, this is my covenant with them," says the LORD. "My Spirit, who is on you, and my words that I have put in your mouth will not depart from your mouth, or from the mouths of your children, or from the mouths of their descendants from this time on and forever," says the LORD.
ISA|60|1|"Arise, shine, for your light has come, and the glory of the LORD rises upon you.
ISA|60|2|See, darkness covers the earth and thick darkness is over the peoples, but the LORD rises upon you and his glory appears over you.
ISA|60|3|Nations will come to your light, and kings to the brightness of your dawn.
ISA|60|4|"Lift up your eyes and look about you: All assemble and come to you; your sons come from afar, and your daughters are carried on the arm.
ISA|60|5|Then you will look and be radiant, your heart will throb and swell with joy; the wealth on the seas will be brought to you, to you the riches of the nations will come.
ISA|60|6|Herds of camels will cover your land, young camels of Midian and Ephah. And all from Sheba will come, bearing gold and incense and proclaiming the praise of the LORD.
ISA|60|7|All Kedar's flocks will be gathered to you, the rams of Nebaioth will serve you; they will be accepted as offerings on my altar, and I will adorn my glorious temple.
ISA|60|8|"Who are these that fly along like clouds, like doves to their nests?
ISA|60|9|Surely the islands look to me; in the lead are the ships of Tarshish, bringing your sons from afar, with their silver and gold, to the honor of the LORD your God, the Holy One of Israel, for he has endowed you with splendor.
ISA|60|10|"Foreigners will rebuild your walls, and their kings will serve you. Though in anger I struck you, in favor I will show you compassion.
ISA|60|11|Your gates will always stand open, they will never be shut, day or night, so that men may bring you the wealth of the nations- their kings led in triumphal procession.
ISA|60|12|For the nation or kingdom that will not serve you will perish; it will be utterly ruined.
ISA|60|13|"The glory of Lebanon will come to you, the pine, the fir and the cypress together, to adorn the place of my sanctuary; and I will glorify the place of my feet.
ISA|60|14|The sons of your oppressors will come bowing before you; all who despise you will bow down at your feet and will call you the City of the LORD, Zion of the Holy One of Israel.
ISA|60|15|"Although you have been forsaken and hated, with no one traveling through, I will make you the everlasting pride and the joy of all generations.
ISA|60|16|You will drink the milk of nations and be nursed at royal breasts. Then you will know that I, the LORD, am your Savior, your Redeemer, the Mighty One of Jacob.
ISA|60|17|Instead of bronze I will bring you gold, and silver in place of iron. Instead of wood I will bring you bronze, and iron in place of stones. I will make peace your governor and righteousness your ruler.
ISA|60|18|No longer will violence be heard in your land, nor ruin or destruction within your borders, but you will call your walls Salvation and your gates Praise.
ISA|60|19|The sun will no more be your light by day, nor will the brightness of the moon shine on you, for the LORD will be your everlasting light, and your God will be your glory.
ISA|60|20|Your sun will never set again, and your moon will wane no more; the LORD will be your everlasting light, and your days of sorrow will end.
ISA|60|21|Then will all your people be righteous and they will possess the land forever. They are the shoot I have planted, the work of my hands, for the display of my splendor.
ISA|60|22|The least of you will become a thousand, the smallest a mighty nation. I am the LORD; in its time I will do this swiftly."
ISA|61|1|The Spirit of the Sovereign LORD is on me, because the LORD has anointed me to preach good news to the poor. He has sent me to bind up the brokenhearted, to proclaim freedom for the captives and release from darkness for the prisoners,
ISA|61|2|to proclaim the year of the LORD's favor and the day of vengeance of our God, to comfort all who mourn,
ISA|61|3|and provide for those who grieve in Zion- to bestow on them a crown of beauty instead of ashes, the oil of gladness instead of mourning, and a garment of praise instead of a spirit of despair. They will be called oaks of righteousness, a planting of the LORD for the display of his splendor.
ISA|61|4|They will rebuild the ancient ruins and restore the places long devastated; they will renew the ruined cities that have been devastated for generations.
ISA|61|5|Aliens will shepherd your flocks; foreigners will work your fields and vineyards.
ISA|61|6|And you will be called priests of the LORD, you will be named ministers of our God. You will feed on the wealth of nations, and in their riches you will boast.
ISA|61|7|Instead of their shame my people will receive a double portion, and instead of disgrace they will rejoice in their inheritance; and so they will inherit a double portion in their land, and everlasting joy will be theirs.
ISA|61|8|"For I, the LORD, love justice; I hate robbery and iniquity. In my faithfulness I will reward them and make an everlasting covenant with them.
ISA|61|9|Their descendants will be known among the nations and their offspring among the peoples. All who see them will acknowledge that they are a people the LORD has blessed."
ISA|61|10|I delight greatly in the LORD; my soul rejoices in my God. For he has clothed me with garments of salvation and arrayed me in a robe of righteousness, as a bridegroom adorns his head like a priest, and as a bride adorns herself with her jewels.
ISA|61|11|For as the soil makes the sprout come up and a garden causes seeds to grow, so the Sovereign LORD will make righteousness and praise spring up before all nations.
ISA|62|1|For Zion's sake I will not keep silent, for Jerusalem's sake I will not remain quiet, till her righteousness shines out like the dawn, her salvation like a blazing torch.
ISA|62|2|The nations will see your righteousness, and all kings your glory; you will be called by a new name that the mouth of the LORD will bestow.
ISA|62|3|You will be a crown of splendor in the LORD's hand, a royal diadem in the hand of your God.
ISA|62|4|No longer will they call you Deserted, or name your land Desolate. But you will be called Hephzibah, and your land Beulah; for the LORD will take delight in you, and your land will be married.
ISA|62|5|As a young man marries a maiden, so will your sons marry you; as a bridegroom rejoices over his bride, so will your God rejoice over you.
ISA|62|6|I have posted watchmen on your walls, O Jerusalem; they will never be silent day or night. You who call on the LORD, give yourselves no rest,
ISA|62|7|and give him no rest till he establishes Jerusalem and makes her the praise of the earth.
ISA|62|8|The LORD has sworn by his right hand and by his mighty arm: "Never again will I give your grain as food for your enemies, and never again will foreigners drink the new wine for which you have toiled;
ISA|62|9|but those who harvest it will eat it and praise the LORD, and those who gather the grapes will drink it in the courts of my sanctuary."
ISA|62|10|Pass through, pass through the gates! Prepare the way for the people. Build up, build up the highway! Remove the stones. Raise a banner for the nations.
ISA|62|11|The LORD has made proclamation to the ends of the earth: "Say to the Daughter of Zion, 'See, your Savior comes! See, his reward is with him, and his recompense accompanies him.'"
ISA|62|12|They will be called the Holy People, the Redeemed of the LORD; and you will be called Sought After, the City No Longer Deserted.
ISA|63|1|Who is this coming from Edom, from Bozrah, with his garments stained crimson? Who is this, robed in splendor, striding forward in the greatness of his strength? "It is I, speaking in righteousness, mighty to save."
ISA|63|2|Why are your garments red, like those of one treading the winepress?
ISA|63|3|"I have trodden the winepress alone; from the nations no one was with me. I trampled them in my anger and trod them down in my wrath; their blood spattered my garments, and I stained all my clothing.
ISA|63|4|For the day of vengeance was in my heart, and the year of my redemption has come.
ISA|63|5|I looked, but there was no one to help, I was appalled that no one gave support; so my own arm worked salvation for me, and my own wrath sustained me.
ISA|63|6|I trampled the nations in my anger; in my wrath I made them drunk and poured their blood on the ground."
ISA|63|7|I will tell of the kindnesses of the LORD, the deeds for which he is to be praised, according to all the LORD has done for us- yes, the many good things he has done for the house of Israel, according to his compassion and many kindnesses.
ISA|63|8|He said, "Surely they are my people, sons who will not be false to me"; and so he became their Savior.
ISA|63|9|In all their distress he too was distressed, and the angel of his presence saved them. In his love and mercy he redeemed them; he lifted them up and carried them all the days of old.
ISA|63|10|Yet they rebelled and grieved his Holy Spirit. So he turned and became their enemy and he himself fought against them.
ISA|63|11|Then his people recalled the days of old, the days of Moses and his people- where is he who brought them through the sea, with the shepherd of his flock? Where is he who set his Holy Spirit among them,
ISA|63|12|who sent his glorious arm of power to be at Moses' right hand, who divided the waters before them, to gain for himself everlasting renown,
ISA|63|13|who led them through the depths? Like a horse in open country, they did not stumble;
ISA|63|14|like cattle that go down to the plain, they were given rest by the Spirit of the LORD. This is how you guided your people to make for yourself a glorious name.
ISA|63|15|Look down from heaven and see from your lofty throne, holy and glorious. Where are your zeal and your might? Your tenderness and compassion are withheld from us.
ISA|63|16|But you are our Father, though Abraham does not know us or Israel acknowledge us; you, O LORD, are our Father, our Redeemer from of old is your name.
ISA|63|17|Why, O LORD, do you make us wander from your ways and harden our hearts so we do not revere you? Return for the sake of your servants, the tribes that are your inheritance.
ISA|63|18|For a little while your people possessed your holy place, but now our enemies have trampled down your sanctuary.
ISA|63|19|We are yours from of old; but you have not ruled over them, they have not been called by your name.
ISA|64|1|Oh, that you would rend the heavens and come down, that the mountains would tremble before you!
ISA|64|2|As when fire sets twigs ablaze and causes water to boil, come down to make your name known to your enemies and cause the nations to quake before you!
ISA|64|3|For when you did awesome things that we did not expect, you came down, and the mountains trembled before you.
ISA|64|4|Since ancient times no one has heard, no ear has perceived, no eye has seen any God besides you, who acts on behalf of those who wait for him.
ISA|64|5|You come to the help of those who gladly do right, who remember your ways. But when we continued to sin against them, you were angry. How then can we be saved?
ISA|64|6|All of us have become like one who is unclean, and all our righteous acts are like filthy rags; we all shrivel up like a leaf, and like the wind our sins sweep us away.
ISA|64|7|No one calls on your name or strives to lay hold of you; for you have hidden your face from us and made us waste away because of our sins.
ISA|64|8|Yet, O LORD, you are our Father. We are the clay, you are the potter; we are all the work of your hand.
ISA|64|9|Do not be angry beyond measure, O LORD; do not remember our sins forever. Oh, look upon us, we pray, for we are all your people.
ISA|64|10|Your sacred cities have become a desert; even Zion is a desert, Jerusalem a desolation.
ISA|64|11|Our holy and glorious temple, where our fathers praised you, has been burned with fire, and all that we treasured lies in ruins.
ISA|64|12|After all this, O LORD, will you hold yourself back? Will you keep silent and punish us beyond measure?
ISA|65|1|"I revealed myself to those who did not ask for me; I was found by those who did not seek me. To a nation that did not call on my name, I said, 'Here am I, here am I.'
ISA|65|2|All day long I have held out my hands to an obstinate people, who walk in ways not good, pursuing their own imaginations-
ISA|65|3|a people who continually provoke me to my very face, offering sacrifices in gardens and burning incense on altars of brick;
ISA|65|4|who sit among the graves and spend their nights keeping secret vigil; who eat the flesh of pigs, and whose pots hold broth of unclean meat;
ISA|65|5|who say, 'Keep away; don't come near me, for I am too sacred for you!' Such people are smoke in my nostrils, a fire that keeps burning all day.
ISA|65|6|"See, it stands written before me: I will not keep silent but will pay back in full; I will pay it back into their laps-
ISA|65|7|both your sins and the sins of your fathers," says the LORD. "Because they burned sacrifices on the mountains and defied me on the hills, I will measure into their laps the full payment for their former deeds."
ISA|65|8|This is what the LORD says: "As when juice is still found in a cluster of grapes and men say, 'Don't destroy it, there is yet some good in it,' so will I do in behalf of my servants; I will not destroy them all.
ISA|65|9|I will bring forth descendants from Jacob, and from Judah those who will possess my mountains; my chosen people will inherit them, and there will my servants live.
ISA|65|10|Sharon will become a pasture for flocks, and the Valley of Achor a resting place for herds, for my people who seek me.
ISA|65|11|"But as for you who forsake the LORD and forget my holy mountain, who spread a table for Fortune and fill bowls of mixed wine for Destiny,
ISA|65|12|I will destine you for the sword, and you will all bend down for the slaughter; for I called but you did not answer, I spoke but you did not listen. You did evil in my sight and chose what displeases me."
ISA|65|13|Therefore this is what the Sovereign LORD says: "My servants will eat, but you will go hungry; my servants will drink, but you will go thirsty; my servants will rejoice, but you will be put to shame.
ISA|65|14|My servants will sing out of the joy of their hearts, but you will cry out from anguish of heart and wail in brokenness of spirit.
ISA|65|15|You will leave your name to my chosen ones as a curse; the Sovereign LORD will put you to death, but to his servants he will give another name.
ISA|65|16|Whoever invokes a blessing in the land will do so by the God of truth; he who takes an oath in the land will swear by the God of truth. For the past troubles will be forgotten and hidden from my eyes.
ISA|65|17|"Behold, I will create new heavens and a new earth. The former things will not be remembered, nor will they come to mind.
ISA|65|18|But be glad and rejoice forever in what I will create, for I will create Jerusalem to be a delight and its people a joy.
ISA|65|19|I will rejoice over Jerusalem and take delight in my people; the sound of weeping and of crying will be heard in it no more.
ISA|65|20|"Never again will there be in it an infant who lives but a few days, or an old man who does not live out his years; he who dies at a hundred will be thought a mere youth; he who fails to reach a hundred will be considered accursed.
ISA|65|21|They will build houses and dwell in them; they will plant vineyards and eat their fruit.
ISA|65|22|No longer will they build houses and others live in them, or plant and others eat. For as the days of a tree, so will be the days of my people; my chosen ones will long enjoy the works of their hands.
ISA|65|23|They will not toil in vain or bear children doomed to misfortune; for they will be a people blessed by the LORD, they and their descendants with them.
ISA|65|24|Before they call I will answer; while they are still speaking I will hear.
ISA|65|25|The wolf and the lamb will feed together, and the lion will eat straw like the ox, but dust will be the serpent's food. They will neither harm nor destroy on all my holy mountain," says the LORD.
ISA|66|1|This is what the LORD says: "Heaven is my throne, and the earth is my footstool. Where is the house you will build for me? Where will my resting place be?
ISA|66|2|Has not my hand made all these things, and so they came into being?" declares the LORD. "This is the one I esteem: he who is humble and contrite in spirit, and trembles at my word.
ISA|66|3|But whoever sacrifices a bull is like one who kills a man, and whoever offers a lamb, like one who breaks a dog's neck; whoever makes a grain offering is like one who presents pig's blood, and whoever burns memorial incense, like one who worships an idol. They have chosen their own ways, and their souls delight in their abominations;
ISA|66|4|so I also will choose harsh treatment for them and will bring upon them what they dread. For when I called, no one answered, when I spoke, no one listened. They did evil in my sight and chose what displeases me."
ISA|66|5|Hear the word of the LORD, you who tremble at his word: "Your brothers who hate you, and exclude you because of my name, have said, 'Let the LORD be glorified, that we may see your joy!' Yet they will be put to shame.
ISA|66|6|Hear that uproar from the city, hear that noise from the temple! It is the sound of the LORD repaying his enemies all they deserve.
ISA|66|7|"Before she goes into labor, she gives birth; before the pains come upon her, she delivers a son.
ISA|66|8|Who has ever heard of such a thing? Who has ever seen such things? Can a country be born in a day or a nation be brought forth in a moment? Yet no sooner is Zion in labor than she gives birth to her children.
ISA|66|9|Do I bring to the moment of birth and not give delivery?" says the LORD. "Do I close up the womb when I bring to delivery?" says your God.
ISA|66|10|"Rejoice with Jerusalem and be glad for her, all you who love her; rejoice greatly with her, all you who mourn over her.
ISA|66|11|For you will nurse and be satisfied at her comforting breasts; you will drink deeply and delight in her overflowing abundance."
ISA|66|12|For this is what the LORD says: "I will extend peace to her like a river, and the wealth of nations like a flooding stream; you will nurse and be carried on her arm and dandled on her knees.
ISA|66|13|As a mother comforts her child, so will I comfort you; and you will be comforted over Jerusalem."
ISA|66|14|When you see this, your heart will rejoice and you will flourish like grass; the hand of the LORD will be made known to his servants, but his fury will be shown to his foes.
ISA|66|15|See, the LORD is coming with fire, and his chariots are like a whirlwind; he will bring down his anger with fury, and his rebuke with flames of fire.
ISA|66|16|For with fire and with his sword the LORD will execute judgment upon all men, and many will be those slain by the LORD.
ISA|66|17|"Those who consecrate and purify themselves to go into the gardens, following the one in the midst of those who eat the flesh of pigs and rats and other abominable things-they will meet their end together," declares the LORD.
ISA|66|18|"And I, because of their actions and their imaginations, am about to come and gather all nations and tongues, and they will come and see my glory.
ISA|66|19|"I will set a sign among them, and I will send some of those who survive to the nations-to Tarshish, to the Libyans and Lydians (famous as archers), to Tubal and Greece, and to the distant islands that have not heard of my fame or seen my glory. They will proclaim my glory among the nations.
ISA|66|20|And they will bring all your brothers, from all the nations, to my holy mountain in Jerusalem as an offering to the LORD -on horses, in chariots and wagons, and on mules and camels," says the LORD. "They will bring them, as the Israelites bring their grain offerings, to the temple of the LORD in ceremonially clean vessels.
ISA|66|21|And I will select some of them also to be priests and Levites," says the LORD.
ISA|66|22|"As the new heavens and the new earth that I make will endure before me," declares the LORD, "so will your name and descendants endure.
ISA|66|23|From one New Moon to another and from one Sabbath to another, all mankind will come and bow down before me," says the LORD.
ISA|66|24|"And they will go out and look upon the dead bodies of those who rebelled against me; their worm will not die, nor will their fire be quenched, and they will be loathsome to all mankind."
