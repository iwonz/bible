EXOD|1|1|以色列 的众儿子各带着家眷，和 雅各 一同来到 埃及 ，他们的名字如下：
EXOD|1|2|吕便 、 西缅 、 利未 、 犹大 、
EXOD|1|3|以萨迦 、 西布伦 、 便雅悯 、
EXOD|1|4|但 、 拿弗他利 、 迦得 、 亚设 。
EXOD|1|5|凡从 雅各 生的，共有七十人。那时， 约瑟 已经在 埃及 。
EXOD|1|6|约瑟 和他所有的兄弟，以及那一代的人都死了。
EXOD|1|7|然而， 以色列 人生养众多，繁衍昌盛，极其强盛，遍满了那地。
EXOD|1|8|有一位不认识 约瑟 的新王兴起，统治 埃及 。
EXOD|1|9|他对自己的百姓说：“看哪， 以色列 人的百姓比我们还多，又比我们强盛。
EXOD|1|10|来吧，让我们机巧地待他们，恐怕他们增多起来，将来若有战争，他们就联合我们的仇敌来攻击我们，然后离开这地去了。”
EXOD|1|11|于是 埃及 人派监工管辖他们，用劳役苦待他们。他们为法老建造储货城，就是 比东 和 兰塞 。
EXOD|1|12|可是越苦待他们，他们就越发增多，更加繁衍， 埃及 人就因 以色列 人愁烦。
EXOD|1|13|埃及 人严厉地强迫 以色列 人做工，
EXOD|1|14|使他们因苦工而生活痛苦；无论是和泥，是做砖，是做田间各样的工，一切的工 埃及 人都严厉地对待他们。
EXOD|1|15|埃及 王又对 希伯来 的接生婆，一个名叫 施弗拉 ，另一个名叫 普阿 的说：
EXOD|1|16|“你们为 希伯来 妇人接生，临盆的时候要注意 ，若是男的，就把他杀了，若是女的，就让她活。”
EXOD|1|17|但是接生婆敬畏上帝，不照 埃及 王的吩咐去做，却让男孩活着。
EXOD|1|18|埃及 王召了接生婆来，对她们说：“你们为什么做这事，让男孩活着呢？”
EXOD|1|19|接生婆对法老说：“因为 希伯来 妇人与 埃及 妇人不同； 希伯来 妇人健壮，接生婆还没有到，她们已经生产了。”
EXOD|1|20|上帝恩待接生婆； 以色列 人增多起来，极其强盛。
EXOD|1|21|接生婆因为敬畏上帝，上帝就叫她们成立家室。
EXOD|1|22|法老吩咐他的众百姓说：“把所生的 每一个男孩都丢到 尼罗河 里去，让所有的女孩存活。”
EXOD|2|1|有一个 利未 家的人娶了一个 利未 女子为妻。
EXOD|2|2|那女人怀孕，生了一个儿子，见他俊美，就把他藏了三个月，
EXOD|2|3|后来不能再藏，就取了一个蒲草箱，抹上柏油和树脂，将孩子放在里面，把箱子搁在 尼罗河 边的芦苇中。
EXOD|2|4|孩子的姊姊远远站着，要知道他究竟会怎样。
EXOD|2|5|法老的女儿来到 尼罗河 边洗澡，她的女仆们在河边行走。她看见在芦苇中的箱子，就派一个使女把它拿来。
EXOD|2|6|她打开箱子，看见那孩子。看哪，男孩在哭，她就可怜他，说：“这是 希伯来 人的一个孩子。”
EXOD|2|7|孩子的姊姊对法老的女儿说：“我去叫一个 希伯来 妇人来作奶妈，替你乳养这孩子，好吗？”
EXOD|2|8|法老的女儿对她说：“去吧！”那女孩就去叫了孩子的母亲来。
EXOD|2|9|法老的女儿对她说：“你把这孩子抱去，替我乳养这孩子，我必给你工钱。”那妇人就把孩子接过来，乳养他。
EXOD|2|10|孩子长大了，妇人把他带到法老的女儿那里，就作了她的儿子。她给孩子起名叫 摩西 ，说：“因我把他从水里拉出来。”
EXOD|2|11|过了一段日子， 摩西 长大了，他出去到他同胞那里，看见他们的劳役。他看见一个 埃及 人打他的同胞，一个 希伯来 人。
EXOD|2|12|他左右观看，见没有人，就把 埃及 人打死了，藏在沙土里。
EXOD|2|13|第二天他出去，看哪，有两个 希伯来 人在打架，他就对那凶恶的人说：“你为什么打你同族的人呢？”
EXOD|2|14|那人说：“谁立你作我们的领袖和审判官呢？难道你要杀我，像杀那 埃及 人一样吗？” 摩西 就惧怕，说：“这事一定是让人知道了。”
EXOD|2|15|法老听见这事，就设法要杀 摩西 。于是 摩西 逃走，躲避法老，到了 米甸 地，坐在井旁。
EXOD|2|16|米甸 的祭司有七个女儿；她们来打水，打满了槽，要给父亲的羊群喝水。
EXOD|2|17|有一些牧羊人来，把她们赶走， 摩西 却起来帮助她们，取水给她们的羊群喝。
EXOD|2|18|她们回到父亲 流珥 那里；他说：“今日你们为何这么快就回来了呢？”
EXOD|2|19|她们说：“有一个 埃及 人来救我们脱离牧羊人的手，他甚至打水给我们的羊群喝。”
EXOD|2|20|他对女儿们说：“那人在哪里？你们为什么撇下他呢？去请他来吃饭吧！”
EXOD|2|21|摩西 愿意和那人同住， 那人就把女儿 西坡拉 给 摩西 为妻。
EXOD|2|22|西坡拉 生了一个儿子， 摩西 给他起名叫 革舜 ，因他说：“我在外地作了寄居者。”
EXOD|2|23|过了许多年， 埃及 王死了。 以色列 人因做苦工，就叹息哀求；他们因苦工所发出的哀声达于上帝。
EXOD|2|24|上帝听见他们的哀声，就记念他与 亚伯拉罕 、 以撒 、 雅各 所立的约。
EXOD|2|25|上帝看顾 以色列 人，上帝是知道的 。
EXOD|3|1|摩西 牧放他岳父 米甸 祭司 叶特罗 的羊群，他领羊群往旷野的那一边去，到了上帝的山，就是 何烈山 。
EXOD|3|2|耶和华的使者在荆棘的火焰中向他显现。 摩西 观看，看哪，荆棘在火中焚烧，却没有烧毁。
EXOD|3|3|摩西 说：“我要转过去看这大异象，这荆棘为何没有烧毁呢？”
EXOD|3|4|耶和华见 摩西 转过去看，上帝就从荆棘里呼叫他说：“ 摩西 ！ 摩西 ！”他说：“我在这里。”
EXOD|3|5|上帝说：“不要靠近这里。把你脚上的鞋脱下来，因为你所站的地方是圣地”。
EXOD|3|6|他又说：“我是你父亲的上帝，是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。” 摩西 蒙上脸，因为怕看上帝。
EXOD|3|7|耶和华说：“我确实看见了我百姓在 埃及 所受的困苦，我也听见了他们因受监工苦待所发的哀声；我确实知道他们的痛苦。
EXOD|3|8|我下来是要救他们脱离 埃及 人的手，领他们从那地上来，到美好与宽阔之地，到流奶与蜜之地，就是 迦南 人、 赫 人、 亚摩利 人、 比利洗 人、 希未 人、 耶布斯 人之地。
EXOD|3|9|现在，看哪， 以色列 人的哀声达到我这里，我也看见 埃及 人怎样欺压他们。
EXOD|3|10|现在，你去，我要差派你到法老那里，把我的百姓 以色列 人从 埃及 领出来。”
EXOD|3|11|摩西 对上帝说：“我是什么人，竟能去见法老，把 以色列 人从 埃及 领出来呢？”
EXOD|3|12|上帝说：“我必与你同在。这就是我差派你去，给你的凭据：你把百姓从 埃及 领出来之后，你们必在这山上事奉上帝。”
EXOD|3|13|摩西 对上帝说：“看哪，我到 以色列 人那里，对他们说：‘你们祖宗的上帝差派我到你们这里来。’他们若对我说：‘他叫什么名字？’我要对他们说什么呢？”
EXOD|3|14|上帝对 摩西 说：“我是自有永有的”；又说：“你要对 以色列 人这样说：‘那自有永有的差派我到你们这里来。’”
EXOD|3|15|上帝又对 摩西 说：“你要对 以色列 人这样说：‘耶和华－你们祖宗的上帝，就是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝差派我到你们这里来。’这是我的名，直到永远；这也是我的称号 ，直到万代。
EXOD|3|16|你去召集 以色列 的长老，对他们说：‘耶和华－你们祖宗的上帝，就是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝向我显现，说：我实在眷顾了你们，眷顾你们在 埃及 的遭遇。
EXOD|3|17|我也曾说：要把你们从 埃及 的困苦中领出来，往 迦南 人、 赫 人、 亚摩利 人、 比利洗 人、 希未 人、 耶布斯 人的地去，就是到流奶与蜜之地。’
EXOD|3|18|他们必听你的话。你和 以色列 的长老要到 埃及 王那里，对他说：‘耶和华－ 希伯来 人的上帝向我们显现，现在求你让我们往旷野去，走三天的路程，为要向耶和华我们的上帝献祭。’
EXOD|3|19|我知道若不用大能的手， 埃及 王不会放你们走。
EXOD|3|20|因此，我必伸出我的手，在 埃及 施行我一切的神迹，击打这地，然后，他才放你们走。
EXOD|3|21|我必使 埃及 人看得起你们，你们离开的时候就不至于空手而去。
EXOD|3|22|每一个妇女必向她的邻舍，以及寄居在她家里的女人，索取金器、银器和衣裳，给你们的儿女穿戴。这样你们就掠夺了 埃及 人。”
EXOD|4|1|摩西 回答说：“看哪！他们不会信我，也不会听我的话，因为他们必说：‘耶和华并没有向你显现。’”
EXOD|4|2|耶和华对 摩西 说：“你手里的是什么？”他说：“是杖。”
EXOD|4|3|耶和华说：“把它丢在地上！”他一丢在地上，杖就变成一条蛇； 摩西 逃走避开它。
EXOD|4|4|耶和华对 摩西 说：“伸出手来，拿住它的尾巴─ 摩西 就伸出手，抓住它，它就在 摩西 的手掌中变为杖─
EXOD|4|5|为了要使他们信耶和华他们祖宗的上帝，就是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝，曾向你显现了。”
EXOD|4|6|耶和华又对他说：“把手放进怀里。”他就把手放进怀里。当他把手抽出来，看哪，手竟然长了痲疯 ，像雪一样白。
EXOD|4|7|耶和华说：“把手放回怀里─他就把手放回怀里。当他把手从怀里再抽出来，看哪，手复原了，与全身的肉一样─
EXOD|4|8|倘若他们不信你，也不听第一个神迹的声音，他们会信第二个神迹的声音。
EXOD|4|9|倘若他们不信这两个神迹，不听你的话，你就从 尼罗河 里取些水，倒在干的地上。你从 尼罗河 里所取的水必在干地上变成血。”
EXOD|4|10|摩西 对耶和华说：“主啊，求求你，我并不是一个能言善道的人，以前这样，就是你对仆人说话以后也是这样，因为我是拙口笨舌的。”
EXOD|4|11|耶和华对他说：“谁造人的口呢？谁使人口哑、耳聋、目明、眼瞎呢？岂不是我－耶和华吗？
EXOD|4|12|现在，去吧，我必赐你口才，指教你应当说的。”
EXOD|4|13|摩西 说：“主啊，求求你，你要藉着谁的手，就差派谁去吧！”
EXOD|4|14|耶和华的怒气向 摩西 发作，说：“你不是有一个哥哥 利未 人 亚伦 吗？我知道他是个能言善道的人。看哪，他正出来迎接你。他一见到你，心里就欢喜。
EXOD|4|15|你要跟他说话，把话放在他的口里，我要赐你口才，也要赐他口才，又要教你们做当做的事。
EXOD|4|16|他要替你向百姓说话；他要当你的口，你要当他的上帝。
EXOD|4|17|你手里要拿这杖，用它来行神迹。”
EXOD|4|18|于是， 摩西 回到他岳父 叶特罗 那里，对他说：“请你让我回 埃及 我同胞那里，看他们还在不在。” 叶特罗 对 摩西 说：“平平安安地去吧！”
EXOD|4|19|耶和华在 米甸 对 摩西 说：“你要回 埃及 去，因为那些寻索你命的人都死了。”
EXOD|4|20|摩西 就带着妻子和两个儿子，让他们骑上驴，回 埃及 地去。 摩西 手里拿着上帝的杖。
EXOD|4|21|耶和华对 摩西 说：“你回到 埃及 去的时候，要留意将我交在你手中的一切奇事行在法老面前。但我要任凭他的心刚硬，他必不放百姓走。
EXOD|4|22|你要对法老说：‘耶和华如此说： 以色列 是我的儿子，我的长子。
EXOD|4|23|我对你说过：放我的儿子走，好事奉我。你还是不肯放他走。看哪，我要杀你头生的儿子。’”
EXOD|4|24|在路上住宿的地方，耶和华遇见 摩西 ，想要杀他。
EXOD|4|25|西坡拉 就拿一块火石，割下她儿子的包皮，碰触 摩西 的脚，说：“你真是我血的新郎了。”
EXOD|4|26|这样，耶和华才放了他。那时， 西坡拉 说：“你因割礼就是血的新郎 了”。
EXOD|4|27|耶和华对 亚伦 说：“你往旷野去迎接 摩西 。”他就去，在上帝的山遇见 摩西 ，就亲他。
EXOD|4|28|摩西 将耶和华差派他所说的话和吩咐他所行的神迹都告诉了 亚伦 。
EXOD|4|29|摩西 和 亚伦 就去召集 以色列 的众长老。
EXOD|4|30|亚伦 将耶和华对 摩西 所说的一切话述说了一遍，又在百姓眼前行了那些神迹，
EXOD|4|31|百姓就信了。他们听见耶和华眷顾 以色列 人，鉴察他们的困苦，就低头敬拜。
EXOD|5|1|后来， 摩西 和 亚伦 去对法老说：“耶和华－ 以色列 的上帝这样说：‘放我的百姓走，好让他们在旷野向我守节。’”
EXOD|5|2|法老说：“耶和华是谁，要我听他的话，让 以色列 人去？我不认识耶和华，也不放 以色列 人走！”
EXOD|5|3|他们说：“ 希伯来 人的上帝已向我们显现了。求你让我们往旷野去，走三天的路程，向耶和华我们的上帝献祭，免得他用瘟疫、刀剑攻击我们。”
EXOD|5|4|埃及 王对他们说：“ 摩西 、 亚伦 ！你们为什么叫百姓不做工呢？去，服你们的劳役吧！”
EXOD|5|5|他又说：“看哪，这地的 以色列 人如今这么多，你们竟然叫他们歇下劳役！”
EXOD|5|6|当天，法老吩咐监工和工头说：
EXOD|5|7|“你们不可照以前一样提供草给百姓做砖，要叫他们自己去捡草。
EXOD|5|8|他们平时做砖的数目，你们仍旧向他们要，一点不可减少，因为他们是懒惰的，所以才呼求说：‘让我们去向我们的上帝献祭。’
EXOD|5|9|你们要把更重的工作加在这些人身上，使他们在其中劳碌，不去理会谎言。”
EXOD|5|10|监工和工头出来对百姓说：“法老这样说：‘我不给你们草，
EXOD|5|11|你们自己在哪里能找到草，就往哪里去找吧！但你们的工作一点也不可减少。’”
EXOD|5|12|于是，百姓分散在 埃及 全地，捡碎秸当草用。
EXOD|5|13|监工催逼他们，说：“你们每天要做完一天的工，与先前有草一样。”
EXOD|5|14|法老的监工击打他们所派的 以色列 工头，说：“为什么昨天和今天你们没有按照以前做砖的数目，完成你们的工作呢？”
EXOD|5|15|以色列 人的工头来哀求法老说：“为什么这样待你的仆人呢？
EXOD|5|16|监工不把草给仆人，并且对我们说：‘做砖吧！’看哪，你仆人挨了打，其实是你百姓的错。”
EXOD|5|17|法老却说：“懒惰，你们真是懒惰！所以你们说：‘让我们去向耶和华献祭吧。’
EXOD|5|18|现在，去做工吧！草是不会给你们，砖却要如数交纳。”
EXOD|5|19|以色列 人的工头听见“你们每天做砖的工作一点也不可减少”，就知道惹上祸了。
EXOD|5|20|他们离开法老出来，正遇见 摩西 和 亚伦 站在那里等候他们，
EXOD|5|21|就向他们说：“愿耶和华鉴察你们，施行判断，因为你们使我们在法老和他臣仆面前有了臭名，把刀递在他们手中来杀我们。”
EXOD|5|22|摩西 回到耶和华那里，说：“主啊，你为什么苦待这百姓呢？为什么差派我呢？
EXOD|5|23|自从我到法老那里，奉你的名说话，他就苦待这百姓，你却一点也没有拯救你的百姓。”
EXOD|6|1|耶和华对 摩西 说：“现在你必看见我向法老所行的事，使他因我大能的手放 以色列 人走，因我大能的手把他们赶出他的地。”
EXOD|6|2|上帝吩咐 摩西 ，对他说：“我是耶和华。
EXOD|6|3|我从前向 亚伯拉罕 、 以撒 、 雅各 显现为全能的上帝；至于我的名耶和华，我未曾让他们知道。
EXOD|6|4|我要与他们坚立我的约，要把 迦南 地，他们寄居的地赐给他们。
EXOD|6|5|我听见 以色列 人被 埃及 人奴役的哀声，我就记念我的约。
EXOD|6|6|所以你要对 以色列 人说：‘我是耶和华；我要除去 埃及 人加给你们的劳役，救你们脱离他们的奴役。我要用伸出来的膀臂，藉严厉的惩罚救赎你们。
EXOD|6|7|我要以你们为我的百姓，我也要作你们的上帝。我除去 埃及 人加给你们的劳役，你们就知道我是耶和华你们的上帝。
EXOD|6|8|我起誓应许给 亚伯拉罕 、 以撒 、 雅各 的地，我要领你们进去，将那地赐给你们为业。我是耶和华。’”
EXOD|6|9|摩西 把这话告诉 以色列 人，但是他们因心里愁烦，又因苦工，就不肯听 摩西 的话。
EXOD|6|10|耶和华吩咐 摩西 说：
EXOD|6|11|“你去对 埃及 王法老说，让 以色列 人离开他的地。”
EXOD|6|12|摩西 在耶和华面前说：“看哪， 以色列 人尚且不听我，法老怎么会听我这不会讲话的人呢？”
EXOD|6|13|耶和华吩咐 摩西 和 亚伦 ，命令他们到 以色列 人和 埃及 王法老那里，把 以色列 人从 埃及 地领出来。
EXOD|6|14|以色列 人族长的名字如下： 以色列 长子 吕便 的儿子是 哈诺 、 法路 、 希斯伦 、 迦米 ；这是 吕便 的家族。
EXOD|6|15|西缅 的儿子是 耶母利 、 雅悯 、 阿辖 、 雅斤 、 琐辖 ，和 迦南 女子生的儿子 扫罗 ；这是 西缅 的家族。
EXOD|6|16|以下是 利未 的儿子按着家谱的名字： 革顺 、 哥辖 、 米拉利 。 利未 一生的岁数是一百三十七岁。
EXOD|6|17|革顺 的儿子按着家族是 立尼 、 示每 。
EXOD|6|18|哥辖 的儿子是 暗兰 、 以斯哈 、 希伯伦 、 乌薛 。 哥辖 一生的岁数是一百三十三岁。
EXOD|6|19|米拉利 的儿子是 抹利 和 母示 ；这是 利未 按着家谱的家族。
EXOD|6|20|暗兰 娶了他父亲的妹妹 约基别 为妻，她为他生了 亚伦 和 摩西 。 暗兰 一生的岁数是一百三十七岁。
EXOD|6|21|以斯哈 的儿子是 可拉 、 尼斐 、 细基利 。
EXOD|6|22|乌薛 的儿子是 米沙利 、 以利撒反 、 西提利 。
EXOD|6|23|亚伦 娶了 亚米拿达 的女儿， 拿顺 的妹妹， 以利沙巴 为妻，她为他生了 拿答 、 亚比户 、 以利亚撒 、 以他玛 。
EXOD|6|24|可拉 的儿子是 亚惜 、 以利加拿 、 亚比亚撒 ；这是 可拉 的家族。
EXOD|6|25|亚伦 的儿子 以利亚撒 娶了 普铁 的一个女儿为妻，她为他生了 非尼哈 。这是 利未 人按着家族的族长。
EXOD|6|26|这就是曾听见耶和华说“把 以色列 人按着队伍从 埃及 地领出来”的 亚伦 和 摩西 ，
EXOD|6|27|对 埃及 王法老说要将 以色列 人从 埃及 领出来的，也是这 摩西 和 亚伦 。
EXOD|6|28|当耶和华在 埃及 地对 摩西 说话的时候，
EXOD|6|29|耶和华对 摩西 说：“我是耶和华；我对你所说的一切话，你都要告诉 埃及 王法老。”
EXOD|6|30|摩西 在耶和华面前说：“看哪，我是不会讲话的人，法老怎么会听我呢？”
EXOD|7|1|耶和华对 摩西 说：“我使你在法老面前像上帝一样，你的哥哥 亚伦 是你的代言人 。
EXOD|7|2|凡我所吩咐你的，你都要说。你的哥哥 亚伦 要对法老说，让 以色列 人离开他的地。
EXOD|7|3|我要使法老的心固执，我也要在 埃及 地多行神迹奇事。
EXOD|7|4|法老必不听从你们，因此我要伸手严厉地惩罚 埃及 ，把我的军队，就是我的百姓 以色列 人从 埃及 地领出来。
EXOD|7|5|我伸手攻击 埃及 ，把 以色列 人从他们中间领出来的时候， 埃及 人就知道我是耶和华。”
EXOD|7|6|摩西 和 亚伦 就去做；他们照耶和华吩咐的去做了。
EXOD|7|7|摩西 和 亚伦 与法老说话的时候， 摩西 八十岁， 亚伦 八十三岁。
EXOD|7|8|耶和华对 摩西 和 亚伦 说：
EXOD|7|9|“法老若吩咐你们说：‘你们行一件奇事吧！’你就对 亚伦 说：‘把杖丢在法老面前！杖会变成蛇。’”
EXOD|7|10|摩西 和 亚伦 到法老那里去，照耶和华所吩咐的去做。 亚伦 把杖丢在法老和他臣仆面前，杖就变成蛇。
EXOD|7|11|法老也召了智慧人和行邪术的人来，这些 埃及 术士也用邪术照样做。
EXOD|7|12|他们各人丢下自己的杖，杖就变成蛇；但 亚伦 的杖吞了他们的杖。
EXOD|7|13|法老心里刚硬，不听 摩西 和 亚伦 ，正如耶和华所说的。
EXOD|7|14|耶和华对 摩西 说：“法老心硬，不肯放百姓走。
EXOD|7|15|明天早晨你要到法老那里去，看哪，他出来往水边去，你要到 尼罗河 边去迎见他，手里拿着那根变过蛇的杖。
EXOD|7|16|你要对他说：‘耶和华－ 希伯来 人的上帝差派我到你这里，说：放我的百姓走，到旷野事奉我。看哪，到如今你还是不听。
EXOD|7|17|耶和华如此说：看哪，我要用我手里的杖击打 尼罗河 中的水，水就变成血；这样，你就知道我是耶和华。
EXOD|7|18|河里的鱼必死，河也要发臭， 埃及 人就厌恶喝这河里的水。’”
EXOD|7|19|耶和华对 摩西 说：“你要对 亚伦 说：‘拿你的杖，伸出你的手在 埃及 所有的水上，在他们的江、河、池塘，所有水聚集的地方上，叫水变成血。在 埃及 全地，无论在木器中，石器中，都必有血。’”
EXOD|7|20|摩西 和 亚伦 就照耶和华所吩咐的去做。 亚伦 在法老和他臣仆眼前举杖击打 尼罗河 里的水，河里的水都变成血了。
EXOD|7|21|河里的鱼死了，河也臭了， 埃及 人就不能喝这河里的水； 埃及 遍地都有了血。
EXOD|7|22|但是， 埃及 的术士也用邪术照样做了；法老心里刚硬，不听 摩西 和 亚伦 ，正如耶和华所说的。
EXOD|7|23|法老转身回宫去，并不把这事放在心上。
EXOD|7|24|所有的 埃及 人都沿着 尼罗河 边挖掘，要找水喝，因为他们不能喝河里的水。
EXOD|7|25|耶和华击打 尼罗河 后，过了七天。
EXOD|8|1|耶和华对 摩西 说：“你要到法老那里，对他说：‘耶和华如此说：放我的百姓走，好事奉我。
EXOD|8|2|你若不肯放他们走，看哪，我必以青蛙之灾击打你的疆土。
EXOD|8|3|尼罗河 要滋生青蛙；这青蛙要上来进你的宫殿和你的卧房，上你的床榻，进你臣仆的房屋，上你百姓的身上，进你的炉灶和你的揉面盆。
EXOD|8|4|这些青蛙要跳上你、你百姓和你众臣仆的身上。’”
EXOD|8|5|耶和华对 摩西 说：“你要对 亚伦 说：‘伸出你手里的杖在江、河、池塘上，把青蛙带上 埃及 地来。’”
EXOD|8|6|亚伦 伸手在 埃及 的众水上，青蛙就上来，遮满了 埃及 地。
EXOD|8|7|术士也用他们的邪术照样去做，把青蛙带上 埃及 地。
EXOD|8|8|法老召 摩西 和 亚伦 来，说：“请你们祈求耶和华使这些青蛙离开我和我的百姓，我就让这百姓去向耶和华献祭。”
EXOD|8|9|摩西 对法老说：“悉听尊便，告诉我何时为你、你臣仆和你的百姓祈求，使青蛙被剪除，离开你和你的宫殿，只留在 尼罗河 里。”
EXOD|8|10|他说：“明天。” 摩西 说：“就照你的话吧，为要叫你知道没有像耶和华我们上帝的，
EXOD|8|11|青蛙必会离开你、你宫殿、你臣仆和你的百姓，只留在 尼罗河 里。”
EXOD|8|12|于是 摩西 和 亚伦 离开法老出去。 摩西 为了青蛙的事呼求耶和华，因为他带来青蛙搅扰法老。
EXOD|8|13|耶和华就照 摩西 的请求去做；在屋里、院中、田间的青蛙都死了。
EXOD|8|14|众人把青蛙聚拢成堆，地就发出臭气。
EXOD|8|15|但法老见灾祸舒缓了，就硬着心，不听从他们，正如耶和华所说的。
EXOD|8|16|耶和华对 摩西 说：“你要对 亚伦 说：‘伸出你的杖击打地上的尘土，使尘土在 埃及 全地变成蚊子 。’”
EXOD|8|17|他们就照样做了。 亚伦 伸出他手里的杖，击打地上的尘土，人和牲畜身上就有了蚊子； 埃及 全地的尘土都变成蚊子了。
EXOD|8|18|术士也用邪术要照样产生蚊子，却做不成。于是人和牲畜的身上都有了蚊子。
EXOD|8|19|术士对法老说：“这是上帝的手指。”法老心里刚硬，不听 摩西 和 亚伦 ，正如耶和华所说的。
EXOD|8|20|耶和华对 摩西 说：“你要清早起来，站在法老面前。看哪，法老来到水边，你就对他说：‘耶和华如此说：放我的百姓走，好事奉我。
EXOD|8|21|你若不放我的百姓走，看哪，我要派成群的苍蝇到你、你臣仆和你百姓身上，进你的宫殿； 埃及 人的房屋和他们所住的地都要满了成群的苍蝇。
EXOD|8|22|那一日，我必把我百姓所住的 歌珊 地分别出来，使那里没有成群的苍蝇，好叫你知道我─耶和华是在全地之中。
EXOD|8|23|我要施行救赎，区隔我的百姓和你的百姓。明天必有这神迹。’”
EXOD|8|24|耶和华就这样做了。大群的苍蝇进入法老的宫殿和他臣仆的房屋；在 埃及 全地，地就因这成群的苍蝇毁坏了。
EXOD|8|25|法老召了 摩西 和 亚伦 来，说：“去，在此地向你们的上帝献祭。”
EXOD|8|26|摩西 说：“这样做是不妥的，因为我们要献给耶和华－我们上帝的祭物是 埃及 人所厌恶的；看哪，我们在 埃及 人眼前献他们所厌恶的，他们岂不拿石头打死我们吗？
EXOD|8|27|我们要遵照耶和华－我们上帝所吩咐我们的，往旷野去，走三天路程，向他献祭。”
EXOD|8|28|法老说：“我可以放你们走，在旷野向耶和华－你们的上帝献祭，只是不可走得太远。你们要为我祈祷。”
EXOD|8|29|摩西 说：“看哪，我要从你这里出去祈求耶和华，使成群的苍蝇明天离开法老、法老的臣仆和法老的百姓；法老却不可再欺骗，不让百姓去向耶和华献祭。”
EXOD|8|30|于是 摩西 离开法老，去祈求耶和华。
EXOD|8|31|耶和华就照 摩西 的请求去做，使成群的苍蝇离开法老、他的臣仆和他的百姓，一只也没有留下。
EXOD|8|32|但这一次法老又硬着心，不放百姓走。
EXOD|9|1|耶和华对 摩西 说：“你要到法老那里，对他说：‘耶和华－ 希伯来 人的上帝如此说：放我的百姓走，好事奉我。
EXOD|9|2|你若不肯放他们走，仍要强留他们，
EXOD|9|3|看哪，耶和华的手必以严重的瘟疫加在你田间的牲畜上，就是在马、驴、骆驼、牛群和羊群的身上。
EXOD|9|4|耶和华却要分别 以色列 的牲畜和 埃及 的牲畜，凡属 以色列 人的，一只都不死。’”
EXOD|9|5|耶和华就设定时间，说：“明天耶和华必在此地行这事。”
EXOD|9|6|第二天，耶和华行了这事。 埃及 的牲畜全都死了，只是 以色列 人的牲畜，一只都没有死。
EXOD|9|7|法老派人去，看哪， 以色列 人的牲畜连一只都没有死。可是法老硬着心，不放百姓走。
EXOD|9|8|耶和华对 摩西 和 亚伦 说：“你们从炉里满满捧出炉灰， 摩西 要在法老眼前把它撒在空中。
EXOD|9|9|这灰要在 埃及 全地变成尘土，使 埃及 全地的人和牲畜身上起泡生疮。”
EXOD|9|10|摩西 和 亚伦 取了炉灰，站在法老面前。 摩西 把它撒在空中，人和牲畜的身上就起泡生疮了。
EXOD|9|11|因为这疮，术士在 摩西 面前站立不住，术士和所有 埃及 人的身上都生了疮。
EXOD|9|12|但耶和华任凭法老的心刚硬，不听 摩西 和 亚伦 ，正如耶和华对 摩西 所说的。
EXOD|9|13|耶和华对 摩西 说：“你要清早起来，站在法老面前，对他说：‘耶和华－ 希伯来 人的上帝如此说：放我的百姓走，好事奉我。
EXOD|9|14|因为这一次我要使一切的灾祸临到你自己，你臣仆和你百姓的身上，为要叫你知道在全地没有像我的。
EXOD|9|15|现在，我若伸手用瘟疫攻击你和你的百姓，你就会从地上除灭了。
EXOD|9|16|然而，我让你存活，是为了要使你看见我的大能，并要使我的名传遍全地。
EXOD|9|17|可是你仍然向我的百姓自高自大，不放他们走。
EXOD|9|18|看哪，明天大约这时候，我必使大量的冰雹降下，这是从 埃及 立国直到如今没有出现过的。
EXOD|9|19|现在，你要派人把你的牲畜和你田间一切所有的带去躲避；任何在田间，无论是人是牲畜没有回到屋内的，冰雹必降在他们身上，他们就必死。’”
EXOD|9|20|法老的臣仆中，惧怕耶和华这话的，就让他的奴仆和牲畜逃进屋里。
EXOD|9|21|但那不把耶和华这话放在心上的，就把他的奴仆和牲畜留在田里。
EXOD|9|22|耶和华对 摩西 说：“你向天伸出你的手，使冰雹降在 埃及 全地，降在 埃及 地的人和牲畜身上，以及田间各样菜蔬上。”
EXOD|9|23|摩西 向天伸杖，耶和华就打雷下雹，有火降到地上；耶和华下雹在 埃及 地上。
EXOD|9|24|那时，有雹，也有火在雹中闪烁，极其严重；自从 埃及 立国以来，全地没有像这样的。
EXOD|9|25|在 埃及 全地，冰雹击打田间所有的人和牲畜，击打一切的菜蔬，也打坏了田间一切的树木。
EXOD|9|26|惟独 以色列 人所住的 歌珊 地没有冰雹。
EXOD|9|27|法老差派人去召 摩西 和 亚伦 来，对他们说：“这一次我犯罪了。耶和华是公义的；我和我的百姓是邪恶的。
EXOD|9|28|请你们祈求耶和华，因上帝的雷轰和冰雹已经够了。我要放你们走，你们不用再留下来了。”
EXOD|9|29|摩西 对他说：“我一出城就向耶和华举起双手；雷必止住，也不再有冰雹，叫你知道地是属于耶和华的。
EXOD|9|30|至于你和你的臣仆，我知道你们仍然不敬畏耶和华上帝。”
EXOD|9|31|那时，亚麻和大麦被摧毁了，因为大麦已经吐穗，亚麻也开了花。
EXOD|9|32|只是小麦和粗麦没有被摧毁，因为它们还没有长成。
EXOD|9|33|摩西 离开法老出了城，向耶和华举起双手，雷和雹就止住，雨也不再下在地上了。
EXOD|9|34|法老见雨、雹、雷止住，又再犯罪；他和他的臣仆都硬着心。
EXOD|9|35|法老的心刚硬，不放 以色列 人走，正如耶和华藉着 摩西 所说的。
EXOD|10|1|耶和华对 摩西 说：“你要到法老那里，因我使他硬着心，也使他臣仆硬着心，为要在他们中间 显出我的这些神迹来，
EXOD|10|2|并要叫你将我严厉对付 埃及 的事，和在他们中间所行的神迹，传于儿子和孙子的耳中，好叫你们知道我是耶和华。”
EXOD|10|3|摩西 和 亚伦 就到法老那里，对他说：“耶和华－ 希伯来 人的上帝这样说：‘你在我面前不肯谦卑要到几时呢？放我的百姓走，好事奉我。
EXOD|10|4|你若不肯放我的百姓走，看哪，明天我要使蝗虫进入你的境内，
EXOD|10|5|遮满地面 ，甚至地也看不见了。它们要吃那冰雹后所剩，就是留给你们的；并且要吃那生长在田间的一切树木。
EXOD|10|6|你的宫殿和你众臣仆的房屋，以及一切 埃及 人的房屋，都要被蝗虫占满；你祖宗和你祖宗的祖宗在世以来，直到今日都没有见过。’” 摩西 就转身离开法老出去。
EXOD|10|7|法老的臣仆对法老说：“这家伙成为我们的罗网要到几时呢？让这些人去事奉耶和华－他们的上帝吧！ 埃及 快要灭亡了，你还不知道吗？”
EXOD|10|8|于是 摩西 和 亚伦 被召回来见法老。法老对他们说：“去，事奉耶和华－你们的上帝吧！但要去的是哪些人呢？”
EXOD|10|9|摩西 说：“我们要带着年老的和年少的同去，要带着我们的儿子和女儿，以及我们的羊群牛群一起去，因为我们要向耶和华守节。”
EXOD|10|10|法老对他们说：“愿耶和华与你们同在吧！我若让你们带着你们的孩子同去，看，灾祸就在你们面前 ！
EXOD|10|11|不可都去！你们壮年人去事奉耶和华吧，因为这是你们所求的。”于是法老把他们从自己面前赶出去。
EXOD|10|12|耶和华对 摩西 说：“你向 埃及 地伸出你的手，使蝗虫上到 埃及 地，吃地上冰雹后所剩一切的植物。”
EXOD|10|13|摩西 就向 埃及 地伸杖；整整一昼一夜，耶和华使东风刮在 埃及 地上，到了早晨，东风把蝗虫刮了来。
EXOD|10|14|蝗虫上到 埃及 全地，落在 埃及 全境，非常厉害；蝗虫这么多，是空前绝后的。
EXOD|10|15|蝗虫遮满地面，地上一片黑暗。它们吃尽了地上一切的植物和冰雹过后所剩树上的果子。 埃及 全地，无论是树木，是田间的植物，连一点绿的也没有留下。
EXOD|10|16|于是法老急忙召了 摩西 和 亚伦 来，说：“我得罪了耶和华－你们的上帝，又得罪了你们。
EXOD|10|17|现在求你，就这一次，饶恕我的罪，祈求耶和华－你们的上帝救我脱离这次的死亡。”
EXOD|10|18|摩西 就离开法老，去祈求耶和华。
EXOD|10|19|耶和华转变风向，使强劲的西风吹来，把蝗虫刮起，吹入 红海 ；在 埃及 全境连一只也没有留下。
EXOD|10|20|但耶和华任凭法老的心刚硬，不放 以色列 人走。
EXOD|10|21|耶和华对 摩西 说：“你向天伸出你的手，使黑暗笼罩 埃及 地；这黑暗甚至可以摸得到。”
EXOD|10|22|摩西 向天伸出他的手，浓密的黑暗就笼罩了 埃及 全地三天之久。
EXOD|10|23|三天内，人人彼此看不见，谁也不敢起身离开原地；但所有 以色列 人住的地方却有光。
EXOD|10|24|法老就召 摩西 来，说：“去，事奉耶和华吧！只是你们的羊群牛群要留下来。你们的孩子可以和你们同去。”
EXOD|10|25|摩西 说：“你必须把祭物和燔祭牲交在我们手中，让我们可以向耶和华我们的上帝献祭。
EXOD|10|26|我们的牲畜也要与我们同去，连一蹄也不留下，因为我们要从牲畜中挑选来事奉耶和华－我们的上帝。未到那里之前，我们还不知道要用什么来事奉耶和华。”
EXOD|10|27|但耶和华任凭法老的心刚硬，法老不肯放他们走。
EXOD|10|28|法老对 摩西 说：“离开我去吧！你要小心，不要再见我的面，因为再见我面的那日，你就必死！”
EXOD|10|29|摩西 说：“就照你说的，我也不要再见你的面了！”
EXOD|11|1|耶和华对 摩西 说：“我要再降一个灾祸给法老和 埃及 ，然后他必让你们离开这里。他放你们走的时候，一定会赶你们全都离开这里。
EXOD|11|2|你要传于百姓耳中，叫他们男的女的各向邻舍索取金器银器。”
EXOD|11|3|耶和华使 埃及 人看得起他的百姓 ，并且 摩西 在 埃及 地，在法老臣仆和百姓眼中看为伟大。
EXOD|11|4|摩西 说：“耶和华如此说：‘约到半夜，我必出去走遍 埃及 。
EXOD|11|5|凡在 埃及 地，从坐宝座的法老到推磨 的婢女所生的长子，以及一切头生的牲畜，都必死。
EXOD|11|6|埃及 全地必有大大的哀号，这将是空前绝后的。
EXOD|11|7|至于 以色列 人中，无论是人是牲畜，连狗也不敢向他们吠叫，使你们知道耶和华区别 埃及 和 以色列 。’
EXOD|11|8|你所有的这些臣仆都要下到我这里，向我下拜说：‘请你和跟从你的百姓都离开吧！’然后我才离开。”于是， 摩西 气愤愤地离开法老出去了。
EXOD|11|9|耶和华对 摩西 说：“法老必不听你们，为了要使我在 埃及 地多行奇事。”
EXOD|11|10|摩西 和 亚伦 在法老面前行了这一切奇事，但耶和华任凭法老的心刚硬，不让 以色列 人离开他的地。
EXOD|12|1|耶和华在 埃及 地对 摩西 和 亚伦 说：
EXOD|12|2|“你们要以本月为正月，为一年之首。
EXOD|12|3|你们要吩咐 以色列 全会众说：本月初十，各人要按着家庭 取羔羊，一家一只羔羊。
EXOD|12|4|若一家的人太少，吃不了一只羔羊，就要按照人数和隔壁的邻舍共取一只；你们要按每人的食量来估算羔羊。
EXOD|12|5|你们要从绵羊或山羊中取一只无残疾、一岁的公羔羊，
EXOD|12|6|要把它留到本月十四日；那日黄昏的时候， 以色列 全会众要把羔羊宰了。
EXOD|12|7|他们要取一些血，涂在他们吃羔羊的房屋两边的门框上和门楣上。
EXOD|12|8|当晚要吃羔羊的肉；要用火烤了，与无酵饼和苦菜一起吃。
EXOD|12|9|不可吃生的，或用水煮的，要把羔羊连头带腿和内脏用火烤了吃。
EXOD|12|10|一点也不可留到早晨；若有留到早晨的，要用火烧了。
EXOD|12|11|你们要这样吃羔羊：腰间束带，脚上穿鞋，手中拿杖，快快地吃。这是耶和华的逾越。
EXOD|12|12|因为那夜我要走遍 埃及 地，把 埃及 地一切头生的，无论是人是牲畜，都击杀了；我要对 埃及 所有的神明施行审判。我是耶和华。
EXOD|12|13|这血要在你们所住的房屋上作记号；我一见这血，就逾越你们。我击打 埃及 地的时候，灾殃必不临到你们身上施行毁灭。”
EXOD|12|14|“你们要记念这日，世世代代守这日为耶和华的节日，作为你们永远的定例。
EXOD|12|15|你们要吃无酵饼七日。第一日要把酵从你们各家中除去，因为从第一日到第七日，任何吃有酵之物的，必从 以色列 中剪除。
EXOD|12|16|第一日当有圣会，第七日也当有圣会。在这两日，任何工作都不可做，只能预备各人的食物，这是惟一可做的工作。
EXOD|12|17|你们要守除酵节，因为我在这一日把你们的军队从 埃及 地领出来。所以，你们要世世代代守这日，立为永远的定例。
EXOD|12|18|从正月十四日晚上，直到二十一日晚上，你们要吃无酵饼。
EXOD|12|19|在你们各家中，七日之内不可有酵，因为凡吃有酵之物的，无论是寄居的，是本地的，必从 以色列 的会中剪除。
EXOD|12|20|任何有酵的物，你们都不可吃；在你们一切的住处要吃无酵饼。”
EXOD|12|21|于是， 摩西 召了 以色列 的众长老来，对他们说：“你们要为家人取羔羊，把逾越的羔羊宰了。
EXOD|12|22|要拿一把牛膝草，蘸盆里的血，把盆里的血涂在门楣上和两边的门框上。直到早晨你们谁也不可出自己家里的门。
EXOD|12|23|因为耶和华要走遍 埃及 ，施行击杀，他看见血在门楣上和两边的门框上，耶和华就必逾越那门，不让灭命者进你们的家，施行击杀。
EXOD|12|24|你们要守这命令，作为你们和你们子孙永远的定例。
EXOD|12|25|日后，你们到了耶和华所应许赐给你们的那地，就要守这礼仪。
EXOD|12|26|你们的儿女对你们说：‘这礼仪是什么意思呢？’
EXOD|12|27|你们就说：‘这是献给耶和华逾越节的祭物。当耶和华击杀 埃及 人的时候，他逾越了 以色列 人在 埃及 的房屋，救了我们各家。’”于是百姓低头敬拜。
EXOD|12|28|以色列 人就去做；他们照耶和华吩咐 摩西 和 亚伦 的去做了。
EXOD|12|29|到了半夜，耶和华把 埃及 地所有头生的，就是从坐宝座的法老，到关在牢里的人的长子，以及一切头生的牲畜，尽都杀了。
EXOD|12|30|法老和他众臣仆，以及所有的 埃及 人，都在夜间起来了。在 埃及 有大大的哀号，因为没有一家不死人的。
EXOD|12|31|夜间，法老召了 摩西 和 亚伦 来，说：“起来！你们和 以色列 人，都离开我的百姓出去，照你们所说的，去事奉耶和华吧！
EXOD|12|32|照你们所说的，连羊群牛群也带走，也为我祝福吧！”
EXOD|12|33|埃及 人催促百姓赶快离开那地，因为 埃及 人说：“我们都快死了。”
EXOD|12|34|百姓就拿着没有发酵的生面，把揉面盆包在衣服中，扛在肩上。
EXOD|12|35|以色列 人照 摩西 的话去做，向 埃及 人索取金器、银器和衣裳。
EXOD|12|36|耶和华使 埃及 人看得起他的百姓， 埃及 人就给了他们所要的。他们就掠夺了 埃及 人。
EXOD|12|37|以色列 人从 兰塞 起程，往 疏割 去。除了小孩，步行的男人约有六十万。
EXOD|12|38|又有许多不同族群的人，以及众多的羊群牛群，和他们一同上去。
EXOD|12|39|他们用 埃及 带出来的生面烤成无酵饼。这生面是没有发酵的；因为他们被催促离开 埃及 ，不能耽延，就没有为自己预备食物。
EXOD|12|40|以色列 人住在 埃及 共四百三十年。
EXOD|12|41|正满四百三十年的那一天，耶和华的全军从 埃及 地出来了。
EXOD|12|42|这是向耶和华守的夜，他领他们出 埃及 地；这是 以色列 众人世世代代要向耶和华守的夜。
EXOD|12|43|耶和华对 摩西 和 亚伦 说：“逾越节的条例是这样：外邦人不可吃这羔羊。
EXOD|12|44|但是你们用银子买来，又受过割礼的奴仆可以吃。
EXOD|12|45|寄居的和雇工都不可吃。
EXOD|12|46|应当在一个屋子里吃，不可把肉带到屋外，骨头一根也不可折断。
EXOD|12|47|以色列 全会众都要守这礼仪。
EXOD|12|48|若有外人寄居在你那里，要向耶和华守逾越节，他所有的男子务要先受割礼，然后才可以当他是本地人，容许他守这礼仪。但未受割礼的都不可吃这羔羊。
EXOD|12|49|本地人和寄居在你们中间的外人当守同一个条例。”
EXOD|12|50|以色列 众人就去做，他们照耶和华吩咐 摩西 和 亚伦 的去做了。
EXOD|12|51|正当那日，耶和华将 以色列 人按着他们的队伍从 埃及 地领了出来。
EXOD|13|1|耶和华吩咐 摩西 说：
EXOD|13|2|“头生的要分别为圣归我； 以色列 中凡头生的，无论是人是牲畜，都是我的。”
EXOD|13|3|摩西 对百姓说：“你们要记念从 埃及 为奴之家出来的这日，因为耶和华用大能的手将你们从这地领出来。有酵之物都不可吃。
EXOD|13|4|亚笔月的这一日你们走出来了。
EXOD|13|5|将来耶和华领你进 迦南 人、 赫 人、 亚摩利 人、 希未 人、 耶布斯 人之地，就是他向你祖宗起誓应许给你的那流奶与蜜之地，那时你要在这一个月守这礼仪。
EXOD|13|6|你要吃无酵饼七日，在第七日要向耶和华守节。
EXOD|13|7|这七日之内，要吃无酵饼；在你的全境内不可见有酵之物，也不可见酵母。
EXOD|13|8|当那日，你要告诉你的儿子说：‘这样做是因为耶和华在我出 埃及 的时候为我所做的事。’
EXOD|13|9|这要在你手上作记号，在你额上 作纪念，使耶和华的教导常在你口中，因为耶和华用大能的手将你从 埃及 领出来。
EXOD|13|10|所以你每年要按着日期守这条例。”
EXOD|13|11|“当耶和华照他向你和你祖宗所起的誓将你领进 迦南 人之地，把那地赐给你的时候，
EXOD|13|12|你要将一切头生的献给耶和华；你牲畜中头生的，公的都归耶和华。
EXOD|13|13|然而，凡头生的驴，你要用羔羊赎回；若不赎它，就要打断它的颈项。你儿子中的长子都要赎出来。
EXOD|13|14|日后，你的儿子问你说：‘这是什么意思？’你就说：‘耶和华用大能的手将我们从 埃及 为奴之家领出来。
EXOD|13|15|那时法老固执，不肯放我们走，耶和华就把 埃及 地所有头生的，无论是人是牲畜，都杀了。因此，我把一切头生的公的牲畜献给耶和华为祭，却将所有头生的儿子赎出来。
EXOD|13|16|这要在你手上作记号，在你额上作经匣 ，因为耶和华用大能的手将我们从 埃及 领出来。’”
EXOD|13|17|法老放百姓走的时候， 非利士 人之地的路虽近，上帝却不领他们从那里走，因为上帝说：“恐怕百姓遇见战争就后悔，转回 埃及 去。”
EXOD|13|18|上帝领百姓绕道而行，走旷野的路到 红海 。 以色列 人出 埃及 地，都带着兵器上去 。
EXOD|13|19|摩西 把 约瑟 的骸骨一起带走；因为 约瑟 曾叫 以色列 人郑重地起誓，对他们说：“上帝必定眷顾你们，你们要把我的骸骨从这里一起带上去。”
EXOD|13|20|他们从 疏割 起程，在旷野边上的 以倘 安营。
EXOD|13|21|耶和华走在他们前面，日间用云柱引领他们的路，夜间用火柱照亮他们，使他们日夜都可以行走。
EXOD|13|22|日间的云柱，夜间的火柱，总不离开百姓的面前。
EXOD|14|1|耶和华吩咐 摩西 说：
EXOD|14|2|“你吩咐 以色列 人转回，要在 比．哈希录 前面， 密夺 和海的中间， 巴力．洗分 的前面安营。你们要在对面，靠近海边安营。
EXOD|14|3|以色列 人这样做，法老必说：‘他们在此地迷了路，旷野把他们困住了。’
EXOD|14|4|我要任凭法老的心刚硬，他要追赶他们。我必在法老和他全军身上得荣耀， 埃及 人就知道我是耶和华。”于是 以色列 人照样做了。
EXOD|14|5|有人报告 埃及 王说：“百姓逃跑了！”法老和他的臣仆对百姓改变了心意，说：“我们放 以色列 人走，不再服事我们，我们怎么会做这种事呢？”
EXOD|14|6|法老就预备战车，带领他的军兵同去，
EXOD|14|7|他带了六百辆特选的战车和 埃及 所有的战车，每辆都有军官。
EXOD|14|8|耶和华任凭 埃及 王法老的心刚硬，他就追赶 以色列 人； 以色列 人却抬起头 来出去了。
EXOD|14|9|埃及 人追赶他们，法老一切的马匹、战车、战车长，与军兵就在海边上，靠近 比．哈希录 ，在 巴力．洗分 的前面，在他们安营的地方追上了。
EXOD|14|10|法老逼近的时候， 以色列 人举目，看哪， 埃及 人追来了，就非常惧怕， 以色列 人向耶和华哀求。
EXOD|14|11|他们对 摩西 说：“难道 埃及 没有坟地，你要把我们带来死在旷野吗？你为什么这样待我们，将我们从 埃及 领出来呢？
EXOD|14|12|我们在 埃及 岂没有对你说过，不要搅扰我们，让我们服事 埃及 人吗？因为服事 埃及 人总比死在旷野好。”
EXOD|14|13|摩西 对百姓说：“不要怕，要站稳，看耶和华今天向你们所要施行的拯救，因为你们今天所看见的 埃及 人必永远不再看见了。
EXOD|14|14|耶和华必为你们争战，你们要安静！”
EXOD|14|15|耶和华对 摩西 说：“你为什么向我哀求呢？你吩咐 以色列 人往前走。
EXOD|14|16|你举手向海伸杖，把水分开。 以色列 人要下到海中，走在干地上。
EXOD|14|17|看哪，我要任凭 埃及 人的心刚硬，他们就跟着下去。我要在法老和他的全军、战车、战车长身上得荣耀。
EXOD|14|18|我在法老和他的战车、战车长身上得荣耀的时候， 埃及 人就知道我是耶和华。”
EXOD|14|19|在 以色列 营前行走的上帝的使者移动，走到他们后面；云也从他们的前面移动，站在他们后面。
EXOD|14|20|它来到 埃及 营和 以色列 营的中间：一边有云和黑暗，另一边它照亮夜晚，整夜彼此不得接近。
EXOD|14|21|摩西 向海伸手，耶和华就用强劲的东风，使海水在一夜间退去，海就成了干地；水分开了。
EXOD|14|22|以色列 人下到海中，走在干地上，水在他们左右成了墙壁。
EXOD|14|23|埃及 人追赶他们，法老一切的马匹、战车和战车长都跟着下到海中。
EXOD|14|24|破晓时分，耶和华从云柱、火柱中了望 埃及 的军兵，使 埃及 的军兵混乱。
EXOD|14|25|他使他们的车轮脱落 ，难以前行， 埃及 人说：“我们从 以色列 人面前逃跑吧！因耶和华为他们作战，攻击 埃及 了。”
EXOD|14|26|耶和华对 摩西 说：“你要向海伸手，使水回流到 埃及 人，他们的战车和战车长身上。”
EXOD|14|27|摩西 就向海伸手，到了天亮的时候，海恢复原状。 埃及 人逃避水的时候，耶和华把他们推入海中。
EXOD|14|28|海水回流，淹没了战车和战车长，以及那些跟着 以色列 人下到海中的法老全军，连一个也没有剩下。
EXOD|14|29|以色列 人却在海中走干地，水在他们的左右成了墙壁。
EXOD|14|30|那一日，耶和华拯救 以色列 脱离 埃及 人的手。 以色列 人看见 埃及 人死在海边。
EXOD|14|31|以色列 人看见耶和华向 埃及 人所施展的大能，百姓就敬畏耶和华，并且信服耶和华和他的仆人 摩西 。
EXOD|15|1|那时， 摩西 和 以色列 人向耶和华唱这歌，说： “我要向耶和华歌唱，因他大大得胜， 将马和骑马的投在海中。
EXOD|15|2|耶和华是我的力量，是我的诗歌， 他也成了我的拯救。 这是我的上帝，我要赞美他； 我父亲的上帝，我要尊崇他。
EXOD|15|3|耶和华是战士； 耶和华是他的名。
EXOD|15|4|“法老的战车、军兵，他已抛在海中； 法老精选的军官都沉于 红海 。
EXOD|15|5|深水淹没他们； 他们好像石头坠到深处。
EXOD|15|6|耶和华啊，你的右手施展能力，大显荣耀； 耶和华啊，你的右手摔碎仇敌。
EXOD|15|7|你大发威严，摧毁了你的敌人； 你发出烈怒，吞灭他们如同碎秸。
EXOD|15|8|因你鼻中的气，水就聚成堆， 大水竖立如垒， 海的中心深水凝结。
EXOD|15|9|仇敌说：‘我要追赶，我要追上， 我要分掳物，在他们身上满足我的心愿， 我要拔刀，亲手毁灭他们。’
EXOD|15|10|你用风一吹，海水就淹没他们； 他们像铅沉在大水之中。
EXOD|15|11|“耶和华啊，众神明中，谁能像你？ 谁能像你，至圣至荣， 可颂可畏，施行奇事！
EXOD|15|12|你伸出右手， 地就吞灭他们。
EXOD|15|13|“你以慈爱引领你所救赎的百姓； 你以能力引导他们到你的圣所。
EXOD|15|14|万民听见就战抖； 疼痛抓住 非利士 的居民。
EXOD|15|15|那时， 以东 的族长惊惶， 摩押 的英雄被战兢抓住， 迦南 所有的居民都融化。
EXOD|15|16|惊骇恐惧临到他们； 耶和华啊，因你膀臂的大能， 他们如石头寂静不动， 等候你百姓过去， 等候你所赎的百姓过去。
EXOD|15|17|你要将他们领进去，栽在你产业的山上， 耶和华啊，就是你为自己所造的住处， 主啊，就是你手所建立的圣所。
EXOD|15|18|耶和华必作王，直到永永远远！”
EXOD|15|19|法老的马匹、战车和战车长下到海中，耶和华使海水回流到他们身上； 以色列 人却走在海中的干地上。
EXOD|15|20|那时， 米利暗 女先知， 亚伦 的姊姊，手里拿着铃鼓；众妇女也跟她出去打鼓跳舞。
EXOD|15|21|米利暗 回应他们： “你们要歌颂耶和华，因他大大得胜， 将马和骑马的投在海中。”
EXOD|15|22|摩西 领 以色列 人从 红海 起程，到了 书珥 的旷野，在旷野走了三天，找不到水。
EXOD|15|23|到了 玛拉 ，他们不能喝 玛拉 的水，因为水是苦的；所以那地名叫 玛拉 。
EXOD|15|24|百姓就向 摩西 发怨言，说：“我们喝什么呢？”
EXOD|15|25|摩西 呼求耶和华，耶和华指示他一棵树 。他把树丢在水里，水就变甜了。 耶和华在那里为他们定了律例、典章，在那里考验他们。
EXOD|15|26|他说：“你若留心听从耶和华－你上帝的话，行我眼中看为正的事，侧耳听我的诫令，遵守我一切的律例，我就不将所加于 埃及 人的疾病加在你身上，因为我是医治你的耶和华。”
EXOD|15|27|他们到了 以琳 ，在那里有十二股水泉，七十棵棕树；他们就在那里的水边安营。
EXOD|16|1|以色列 全会众从 以琳 起程，在出 埃及 之后第二个月十五日到了 以琳 和 西奈 中间， 汛 的旷野。
EXOD|16|2|以色列 全会众在旷野向 摩西 和 亚伦 发怨言。
EXOD|16|3|以色列 人对他们说：“我们宁愿在 埃及 地死在耶和华手中！那时我们坐在肉锅旁，吃饼得饱。你们却将我们领出来，到这旷野，要叫这全会众都饿死啊！”
EXOD|16|4|耶和华对 摩西 说：“看哪，我要从天降食物给你们。百姓可以出去，每天收集当天的分量。这样，我就可以考验他们是否遵行我的指示。
EXOD|16|5|到第六天，他们预备食物，所收集的分量要比每天所收的多一倍。”
EXOD|16|6|摩西 和 亚伦 对 以色列 众人说：“到了晚上，你们就知道是耶和华将你们从 埃及 地领出来的。
EXOD|16|7|早晨，你们要看见耶和华的荣耀，因为耶和华听见你们向他所发的怨言了。我们算什么，你们竟然向我们发怨言呢？”
EXOD|16|8|摩西 又说：“耶和华晚上必给你们肉吃，早晨必给你们食物得饱，因为耶和华已经听见你们向他所发的怨言。我们算什么呢？你们的怨言不是向我们发的，而是向耶和华发的。”
EXOD|16|9|摩西 对 亚伦 说：“你对 以色列 全会众说：‘你们来到耶和华面前，因为他已经听见你们的怨言了。’”
EXOD|16|10|亚伦 正对 以色列 全会众说话的时候，他们转向旷野，看哪，耶和华的荣光在云中显现。
EXOD|16|11|耶和华吩咐 摩西 说：
EXOD|16|12|“我已经听见 以色列 人的怨言了。你要对他们说：‘到黄昏的时候 ，你们要吃肉，早晨也必有食物得饱。你们就知道我是耶和华－你们的上帝。’”
EXOD|16|13|到了晚上，有鹌鹑上来，遮满营地；早晨，营地周围有一层露水。
EXOD|16|14|那一层露水蒸发之后，看哪，旷野的表面出现了小圆物，好像地上的薄霜一样。
EXOD|16|15|以色列 人看见了，不知道是什么，就彼此说：“这是什么？ ” 摩西 对他们说：“这是耶和华给你们吃的食物。
EXOD|16|16|耶和华所吩咐的是这样：‘你们每个人要按自己的食量收集，各人要为帐棚里的人收集，按照人口数每个人一俄梅珥。’”
EXOD|16|17|以色列 人就照样去做；有的收多，有的收少。
EXOD|16|18|用俄梅珥量一量，多收的没有余，少收的也没有缺；各人都按着自己的食量收集。
EXOD|16|19|摩西 对他们说：“任何人都不可以把所收的留到早晨。”
EXOD|16|20|然而他们不听从 摩西 ，当中有人把食物留到早晨，食物就生虫发臭了。 摩西 就向他们发怒。
EXOD|16|21|他们每日早晨按着各人的食量收集；太阳一发热，食物就融化了。
EXOD|16|22|到第六天，他们收集了双倍的食物，每个人二俄梅珥。会众的官长来告诉 摩西 ，
EXOD|16|23|摩西 对他们说：“耶和华吩咐：‘明天是安息日，是向耶和华守的圣安息日。你们要烤的就烤，要煮的就煮，所剩下的都留到早晨。’”
EXOD|16|24|他们就照 摩西 的吩咐把剩下的留到早晨，这些食物既不发臭，里头也没有生虫。
EXOD|16|25|摩西 说：“你们今天就吃这些吧！因为今天是向耶和华守的安息日，你们在野外必找不着食物了。
EXOD|16|26|六天可以收集，第七天是安息日，这一天什么也没有了。”
EXOD|16|27|第七天，百姓中有人出去收，什么也找不着。
EXOD|16|28|耶和华对 摩西 说：“你们不肯遵守我的诫令和教导，要到几时呢？
EXOD|16|29|你们看，耶和华既然将安息日赐给你们，所以第六天他就赐给你们两天的食物，第七天各人都要留在自己的地方，不许任何人从这里出去。”
EXOD|16|30|于是百姓在第七天安息了。
EXOD|16|31|以色列 家给这食物取名叫吗哪，它的样子像芫荽子，颜色是白的，吃起来像和蜜的薄饼。
EXOD|16|32|摩西 说：“耶和华所吩咐的是这样：‘要装满一俄梅珥的吗哪留给你们的后代，使他们可以看见我领你们出 埃及 地的时候，在旷野所给你们吃的食物。’”
EXOD|16|33|摩西 对 亚伦 说：“你拿一个罐子，装满一俄梅珥的吗哪，存在耶和华面前，留给你们的后代。”
EXOD|16|34|耶和华怎么吩咐 摩西 ， 亚伦 就照样做，把吗哪存留作见证 。
EXOD|16|35|以色列 人吃吗哪共四十年，直到进入有人居住的地方；他们吃吗哪，直到 迦南 地的边境。
EXOD|16|36|一俄梅珥是一伊法的十分之一。
EXOD|17|1|以色列 全会众遵照耶和华的吩咐，从 汛 的旷野一段一段地往前行。他们在 利非订 安营，但百姓没有水喝。
EXOD|17|2|百姓就与 摩西 争闹，说：“给我们水喝吧！” 摩西 对他们说：“你们为什么与我争闹呢？你们为什么试探耶和华呢？”
EXOD|17|3|百姓在那里口渴要喝水，就向 摩西 发怨言，说：“你为什么把我们从 埃及 领出来，使我们和我们的儿女，以及牲畜都渴死呢？”
EXOD|17|4|摩西 就呼求耶和华说：“我要怎样对待这百姓呢？他们差一点就要拿石头打死我了。”
EXOD|17|5|耶和华对 摩西 说：“你带着 以色列 的几个长老，走在百姓前面，手里拿着你先前击打 尼罗河 的杖，去吧！
EXOD|17|6|看哪，我要在 何烈 的磐石那里，站在你面前。你要击打磐石，水就会从磐石流出来，给百姓喝。” 摩西 就在 以色列 的长老眼前这样做了。
EXOD|17|7|他给那地方起名叫 玛撒 ，又叫 米利巴 ，因为 以色列 人在那里争闹，并且试探耶和华，说：“耶和华是否在我们中间呢？”
EXOD|17|8|那时， 亚玛力 来到 利非订 ，和 以色列 争战。
EXOD|17|9|摩西 对 约书亚 说：“你为我们选出人来，出去和 亚玛力 争战。明天我要站在山顶上，手里拿着上帝的杖。”
EXOD|17|10|于是， 约书亚 照着 摩西 对他所说的话去做，和 亚玛力 争战。 摩西 、 亚伦 和 户珥 都上了山顶。
EXOD|17|11|摩西 何时举手， 以色列 就得胜；何时垂手， 亚玛力 就得胜。
EXOD|17|12|但 摩西 的双手沉重，他们就搬一块石头来放在他下面，他就坐在上面。 亚伦 与 户珥 扶着他的手，一个在这边，一个在那边，他的手就稳住，直到日落。
EXOD|17|13|约书亚 用刀打败了 亚玛力 和他的百姓。
EXOD|17|14|耶和华对 摩西 说：“你要把这事记录在书上作纪念，又念给 约书亚 听：我要把 亚玛力 的名字从天下全然涂去。”
EXOD|17|15|摩西 筑了一座坛，起名叫“耶和华尼西 ”。
EXOD|17|16|他说：“我指着耶和华的宝座发誓 ，耶和华必世世代代和 亚玛力 争战。”
EXOD|18|1|摩西 的岳父， 米甸 祭司 叶特罗 ，听见上帝为 摩西 和为他百姓 以色列 所行的一切事，就是耶和华将 以色列 从 埃及 领了出来。
EXOD|18|2|摩西 的岳父 叶特罗 带着 西坡拉 ，就是 摩西 先前送回家的妻子，
EXOD|18|3|又带着她的两个儿子：一个名叫 革舜 ，因为 摩西 说：“我在外地作了寄居者”；
EXOD|18|4|另一个名叫 以利以谢 ，因为他说：“我父亲的上帝帮助我，救我脱离法老的刀。”
EXOD|18|5|摩西 的岳父 叶特罗 带着 摩西 的妻子和两个儿子来到上帝的山，就是 摩西 在旷野安营的地方。
EXOD|18|6|他对 摩西 说：“我是 你岳父 叶特罗 ，带着你的妻子和两个儿子来到你这里。”
EXOD|18|7|摩西 迎接他的岳父，向他下拜，亲他，彼此问安，然后进入帐棚。
EXOD|18|8|摩西 将耶和华为 以色列 的缘故向法老和 埃及 人所行的一切事，他们在路上遭遇的一切艰难，以及耶和华怎样搭救他们，都述说给他的岳父听。
EXOD|18|9|叶特罗 因耶和华待 以色列 的一切恩惠，就是拯救他们脱离 埃及 人的手，就非常喜乐。
EXOD|18|10|叶特罗 说：“耶和华是应当称颂的，他救了你们脱离 埃及 人和法老的手，将这百姓从 埃及 人的手里救出来 。
EXOD|18|11|现在，从 埃及 人狂傲地对待 以色列 人这件事上，我知道耶和华比万神更大。”
EXOD|18|12|摩西 的岳父 叶特罗 把燔祭和祭物献给上帝。 亚伦 和 以色列 的众长老都来了，与 摩西 的岳父在上帝面前吃饭。
EXOD|18|13|第二天， 摩西 坐着审判百姓，百姓从早到晚站在 摩西 的旁边。
EXOD|18|14|摩西 的岳父看见他为百姓所做的一切事，就说：“你为百姓所做的，这是什么事呢？你为什么独自一人坐着，而众百姓从早到晚都站在你旁边呢？”
EXOD|18|15|摩西 对岳父说：“这是因为百姓到我这里来求问上帝。
EXOD|18|16|他们有事的时候，就到我这里来，我就在双方之间作判决；我又叫他们知道上帝的律例和法度。”
EXOD|18|17|摩西 的岳父对他说：“你这样做不好。
EXOD|18|18|你和这些与你在一起的百姓都必疲惫，因为这事太重，你独自一人做不了。
EXOD|18|19|现在，听我的话，我给你出个主意，愿上帝与你同在。你要代替百姓到上帝面前，将事件带到上帝那里，
EXOD|18|20|又要用律例和法度警戒他们，指示他们当行的道，当做的事。
EXOD|18|21|你也要从百姓中选出有才能的人，敬畏上帝、诚实可靠、恨恶不义之财的人，派他们作千夫长、百夫长、五十夫长、十夫长来管理百姓。
EXOD|18|22|他们要随时审判百姓；重大的事要送到你这里，小事就由他们自行判决。这样，你就可以轻省一些，他们可以与你分担。
EXOD|18|23|你若这样做，上帝也这样吩咐你，你就能承受得住，众百姓也可以和睦地回到自己的地方。”
EXOD|18|24|摩西 听了他岳父的话，照着他所说的一切去做。
EXOD|18|25|摩西 从 以色列 人中选出有才能的人，立他们为百姓的领袖，作千夫长、百夫长、五十夫长、十夫长。
EXOD|18|26|他们随时审判百姓：难断的事就送到 摩西 那里，各样小事就由他们自行判决。
EXOD|18|27|于是， 摩西 给他的岳父送行，他就回到本地去了。
EXOD|19|1|以色列 人出 埃及 地以后，第三个月的初一，就在那一天他们来到了 西奈 的旷野。
EXOD|19|2|他们从 利非订 起程，来到 西奈 的旷野，在那里的山下安营。
EXOD|19|3|摩西 到上帝那里，耶和华从山上呼唤他说：“你要这样告诉 雅各 家，对 以色列 人说：
EXOD|19|4|‘我向 埃及 人所行的事，你们都看见了， 我如鹰将你们背在翅膀上，带你们来归我。
EXOD|19|5|如今你们若真的听从我的话，遵守我的约，就要在万民中作属我的子民 ，因为全地都是我的。
EXOD|19|6|你们要归我作祭司的国度，为神圣的国民。’这些话你要告诉 以色列 人。”
EXOD|19|7|摩西 去召了百姓中的长老来，将耶和华吩咐他的话当面告诉他们。
EXOD|19|8|百姓都同声回答：“凡耶和华所说的，我们一定遵行。” 摩西 就将百姓的话回覆耶和华。
EXOD|19|9|耶和华对 摩西 说：“看哪，我要在密云中临到你那里，叫百姓在我与你说话的时候可以听见，就可以永远相信你了。”于是， 摩西 将百姓的话禀告耶和华。
EXOD|19|10|耶和华对 摩西 说：“你往百姓那里去，使他们今天明天分别为圣，又叫他们洗衣服。
EXOD|19|11|第三天要预备好，因为第三天耶和华要在众百姓眼前降临在 西奈山 。
EXOD|19|12|你要在山的周围给百姓划定界限，说：‘你们当谨慎，不可上山去，也不可摸山的边界。凡摸这山的，必被处死。
EXOD|19|13|不可用手碰他，要用石头打死，或射死；无论是人是牲畜，都不可活。’到角声拉长的时候，他们才可到山脚来。”
EXOD|19|14|摩西 下山到百姓那里去，使他们分别为圣，他们就洗衣服。
EXOD|19|15|他对百姓说：“第三天要预备好；不可亲近女人。”
EXOD|19|16|到了第三天早晨，山上有雷轰、闪电和密云，并且角声非常响亮，营中的百姓尽都战抖。
EXOD|19|17|摩西 率领百姓出营迎见上帝，都站在山下。
EXOD|19|18|西奈山 全山冒烟，因为耶和华在火中降临山上。山的烟雾上腾，仿佛烧窑，整座山剧烈震动。
EXOD|19|19|角声越来越响， 摩西 说话，上帝以声音回答他。
EXOD|19|20|耶和华降临在 西奈山 顶上，耶和华召 摩西 上山顶， 摩西 就上去了。
EXOD|19|21|耶和华对 摩西 说：“你下去警告百姓，免得他们闯过来看耶和华，就会有许多人死亡。
EXOD|19|22|那些亲近耶和华的祭司也要把自己分别为圣，免得耶和华忽然出来击杀他们。”
EXOD|19|23|摩西 对耶和华说：“百姓不能上 西奈山 ，因为你已经警告我们说：‘要在山的周围划定界限，使山成圣。’”
EXOD|19|24|耶和华对他说：“下去吧，你要和 亚伦 一起上来；只是祭司和百姓不可闯上来到耶和华这里，免得耶和华忽然出来击杀他们。”
EXOD|19|25|于是， 摩西 下到百姓那里告诉他们。
EXOD|20|1|上帝吩咐这一切的话，说：
EXOD|20|2|“我是耶和华－你的上帝，曾将你从 埃及 地为奴之家领出来。
EXOD|20|3|“除了我以外，你不可有别的神。
EXOD|20|4|“不可为自己雕刻偶像，也不可做什么形像，仿佛上天、下地和地底下水中的百物。
EXOD|20|5|不可跪拜那些像，也不可事奉它们，因为我耶和华─你的上帝是忌邪 的上帝。恨我的，我必惩罚他们的罪，自父及子，直到三、四代；
EXOD|20|6|爱我，守我诫命的，我必向他们施慈爱，直到千代。
EXOD|20|7|“不可妄称耶和华－你上帝的名，因为妄称耶和华名的，耶和华必不以他为无罪。
EXOD|20|8|“当记念安息日，守为圣日。
EXOD|20|9|六日要劳碌做你一切的工，
EXOD|20|10|但第七日是向耶和华─你的上帝当守的安息日。这一日你和你的儿女、奴仆、婢女、牲畜，以及你城里寄居的客旅，都不可做任何的工。
EXOD|20|11|因为六日之内，耶和华造天、地、海和其中的万物，第七日就安息了；所以耶和华赐福与安息日，定为圣日。
EXOD|20|12|“当孝敬父母，使你的日子在耶和华－你上帝所赐你的地上得以长久。
EXOD|20|13|“不可杀人。
EXOD|20|14|“不可奸淫。
EXOD|20|15|“不可偷盗。
EXOD|20|16|“不可做假见证陷害你的邻舍。
EXOD|20|17|“不可贪恋你邻舍的房屋；不可贪恋你邻舍的妻子、奴仆、婢女、牛驴，以及他一切所有的。”
EXOD|20|18|众百姓见雷轰、闪电、角声、山上冒烟，百姓看见 就都战抖，远远站着。
EXOD|20|19|他们对 摩西 说：“请你向我们说话，我们必听；不要让上帝向我们说话，免得我们死亡。”
EXOD|20|20|摩西 对百姓说：“不要害怕；因为上帝降临是要考验你们，要你们敬畏他，不致犯罪。”
EXOD|20|21|于是百姓远远站着，但 摩西 却挨近上帝所在的幽暗中。
EXOD|20|22|耶和华对 摩西 说：“你要向 以色列 人这样说：‘你们亲自看见我从天上向你们说话了。
EXOD|20|23|你们不可为我制造偶像，不可为自己造任何金银的神像。
EXOD|20|24|你要为我筑一座土坛，在上面献牛羊为燔祭和平安祭。凡在我叫你记念我名的地方，我必到那里赐福给你。
EXOD|20|25|你若为我筑一座石坛，不可用凿过的石头，因为你在石头上动了工具，就使坛污秽了。
EXOD|20|26|你不可用台阶上我的坛，免得露出你的下体来。’”
EXOD|21|1|“你在百姓面前所要立的典章是这样：
EXOD|21|2|“你若买 希伯来 人作奴仆，他服事你六年，第七年他可以自由，白白地离去。
EXOD|21|3|他若单身来就可以单身去；他若是有妻子的，他的妻子可以同他离去。
EXOD|21|4|若他主人给他娶了妻，妻子为他生了儿子或女儿，妻子和儿女要归主人，他要独自离去。
EXOD|21|5|倘若奴仆声明：‘我爱我的主人和我的妻子儿女，不愿意自由离去。’
EXOD|21|6|他的主人就要带他到审判官 前，再带他到门或门框那里，用锥子穿他的耳朵，他就要永远服事主人。
EXOD|21|7|“人若卖女儿作婢女，婢女不可像男的奴仆那样离去。
EXOD|21|8|主人若选定她归自己，后来看不顺眼，就要允许她赎身；主人既然对她失信，就没有权柄把她卖给外邦人。
EXOD|21|9|主人若选定她给自己的儿子，就当照女儿的规矩对待她。
EXOD|21|10|若另娶一个，她的饮食、衣服和房事不可减少。
EXOD|21|11|若不向她行这三样，她就可以白白离去，不必付赎金。”
EXOD|21|12|“打人致死的，必被处死。
EXOD|21|13|他若不是出于预谋 ，而是上帝交在他手中，我就设立一个地方，让他可以逃到那里。
EXOD|21|14|人若蓄意用诡计杀了他的邻舍，就是逃到我的坛那里，也当把他捉去处死。
EXOD|21|15|“打父母的，必被处死。
EXOD|21|16|“诱拐人口的，无论是把人卖了，或是扣留在他手中，必被处死。
EXOD|21|17|“咒骂父母的，必被处死。
EXOD|21|18|“人若彼此争吵，一个用石头或拳头打另一个，被打的人没有死去，却要躺卧在床，
EXOD|21|19|若他还能起来扶杖行走，那打他的可免处刑，却要赔偿他不能工作的损失，并要把他完全医好。
EXOD|21|20|“人若用棍子打奴仆或婢女，当场死在他的手下，他必受报应。
EXOD|21|21|若能撑过一两天，主人就不必受惩罚，因为那是他的财产。
EXOD|21|22|“人若彼此打斗，伤害有孕的妇人，以致胎儿掉了出来，随后却无别的伤害，那伤害她的人，总要按妇人的丈夫所提出的，照审判官所裁定的赔偿。
EXOD|21|23|若有别的伤害，就要以命抵命，
EXOD|21|24|以眼还眼，以牙还牙，以手还手，以脚还脚，
EXOD|21|25|以灼伤还灼伤，以损伤还损伤，以鞭打还鞭打。
EXOD|21|26|“人若打奴仆或婢女的眼睛，毁了一只，就要因他的眼让他自由离去。
EXOD|21|27|若打掉了奴仆或婢女的一颗牙，就要因他的牙让他自由离去。”
EXOD|21|28|“牛若抵死男人或女人，总要用石头打死那牛，却不可吃它的肉；牛的主人可免处刑。
EXOD|21|29|倘若那牛向来是抵人的，牛的主人虽然受过警告，仍不把它拴好，以致把男人或女人抵死，牛要用石头打死，主人也要被处死。
EXOD|21|30|若罚他付赎命的赔款，他就要照所罚的数目赎他的命。
EXOD|21|31|牛若抵了男孩或女孩，也要照这条例处理。
EXOD|21|32|牛若抵了奴仆或婢女，就要把三十舍客勒银子给他的主人，牛要用石头打死。
EXOD|21|33|“人若敞开井口，或挖井不盖住它，有牛或驴掉进井里，
EXOD|21|34|井的主人要拿钱赔偿牲畜的主人，死牲畜要归自己。
EXOD|21|35|“人的牛若抵死邻舍的牛，他们就要卖了那活牛，平分价钱；也要平分死牛。
EXOD|21|36|若这牛向来是以好抵人出名的，主人竟不把牛拴好，他必要以牛赔牛，死牛却归自己。”
EXOD|22|1|“人若偷牛或羊，无论是宰了或卖了，他就要以五牛赔一牛， 四羊赔一羊。
EXOD|22|2|贼挖洞，若被发现而被打死，打的人没有流血的罪。
EXOD|22|3|若太阳已经出来，打的人就有流血的罪。贼总要赔偿，若他一无所有，就要被卖来还他所偷的东西。
EXOD|22|4|若发现他所偷的，无论是牛、驴，或羊，在他手中还活着，他就要加倍赔偿。
EXOD|22|5|“人若在田间或葡萄园里牧放牲畜，任凭牲畜上别人田里去吃 ，他就要拿自己田间和葡萄园里上好的赔偿。
EXOD|22|6|“若火冒出，延烧到荆棘，以致将堆积的禾捆，直立的庄稼，或田地，都烧尽了，那点火的必要赔偿。
EXOD|22|7|“人若将银钱或物件托邻舍保管，东西从这人的家中被偷去，若找到了贼，贼要加倍赔偿；
EXOD|22|8|若找不到贼，这家的主人就要到审判官 那里，声明 自己没有伸手拿邻舍的物件。
EXOD|22|9|“关于任何侵害的案件，无论是为牛、驴、羊、衣服，或任何失物，有一人说：‘这是我的’，双方就要将案件带到审判官面前，审判官定谁有罪，谁就要加倍赔偿给他的邻舍。
EXOD|22|10|“人将驴、牛、羊，或别的牲畜托邻舍看管，若牲畜死亡，受了伤，或被抢走，无人看见，
EXOD|22|11|双方要在耶和华前起誓，受托人要表明自己没有伸手拿邻舍的东西，原主要接受誓言，受托人不必赔偿。
EXOD|22|12|牲畜若从受托人那里被偷去，他就要赔偿原主；
EXOD|22|13|若被野兽撕碎，受托人要带回来作证据，被撕碎的就不必赔偿。
EXOD|22|14|“人若向邻舍借牲畜 ，所借的或伤或死，原主没有在场，借的人总要赔偿。
EXOD|22|15|若原主在场，借的人不必赔偿；若是租用的，只要付租金 。”
EXOD|22|16|“人若引诱没有订婚的处女，与她同寝，他就必须交出聘礼，娶她为妻。
EXOD|22|17|若女子的父亲坚决不将女子给他，他就要按着处女的聘礼交出钱来。
EXOD|22|18|“行邪术的女人，不可让她存活。
EXOD|22|19|“凡与兽交合的，必被处死。
EXOD|22|20|“向别神献祭，不单单献给耶和华的，那人必要灭绝。
EXOD|22|21|“不可亏待寄居的，也不可欺压他，因为你们在 埃及 地也作过寄居的。
EXOD|22|22|不可苛待寡妇和孤儿；
EXOD|22|23|若你确实苛待他，他向我苦苦哀求，我一定会听他的呼求，
EXOD|22|24|并要发烈怒，用刀杀你们，使你们的妻子成为寡妇，儿女成为孤儿。
EXOD|22|25|“我的子民中有困苦人在你那里，你若借钱给他，不可如放债的向他取利息。
EXOD|22|26|你果真拿了邻舍的外衣作抵押，也要在日落前还给他；
EXOD|22|27|因为他只有这一件用来作被子，是他蔽体的衣服。他还可以拿什么睡觉呢？当他哀求我，我就应允，因为我是有恩惠的。
EXOD|22|28|“不可毁谤上帝；也不可诅咒你百姓的领袖。
EXOD|22|29|“不可迟延献你的庄稼、酒和油 。 “要将你头生的儿子归给我。
EXOD|22|30|你的牛羊也要照样做：七天当跟着它母亲，第八天你要把它归给我。
EXOD|22|31|“你们要分别为圣归给我。因此，田间被野兽撕裂的肉，你们不可吃，要把它丢给狗。”
EXOD|23|1|“不可散布谣言；不可与恶人连手作恶意的见证。
EXOD|23|2|不可附和群众作恶；不可在诉讼中附和群众歪曲公正，作歪曲的见证；
EXOD|23|3|也不可在诉讼中偏袒贫寒人。
EXOD|23|4|“若遇见你仇敌的牛或驴迷了路，务必牵回来交给他。
EXOD|23|5|若看见恨你的人的驴被压在重驮之下，不可走开，务要和他一同卸下驴的重驮。
EXOD|23|6|“不可在贫穷人的诉讼中屈枉正直。
EXOD|23|7|当远离诬告的事。不可杀害无辜和义人，因我必不以恶人为义。
EXOD|23|8|不可接受贿赂，因为贿赂能使明眼人变瞎，又能曲解义人的证词。
EXOD|23|9|“不可欺压寄居的，因为你们在 埃及 地作过寄居的，知道寄居者的心情。”
EXOD|23|10|“六年你要耕种田地，收集地的出产。
EXOD|23|11|只是第七年你要让地歇息，不耕不种，使你百姓中的贫穷人有吃的；他们吃剩的，野兽可以吃。你的葡萄园和橄榄园也要照样办理。
EXOD|23|12|“六日你要做工，第七日要安息，使牛、驴可以歇息，也让你使女的儿子和寄居的可以恢复精力。
EXOD|23|13|“凡我对你们说的话，你们都要谨守。别神的名，你不可提，也不可用口说给人听。”
EXOD|23|14|“一年三次，你要向我守节。
EXOD|23|15|你要守除酵节，照我所吩咐你的，在亚笔月内所定的日期吃无酵饼七天，因为你是在这月离开了 埃及 。谁也不可空手来朝见我。
EXOD|23|16|你要守收割节，收田间所种、劳碌所得初熟之物。你年底收藏田间劳碌所得时，要守收藏节。
EXOD|23|17|所有的男丁都要一年三次朝见主耶和华。
EXOD|23|18|“不可将我祭牲的血和有酵之物一同献上，也不可将我节期中祭牲的脂肪留到早晨。
EXOD|23|19|“要把地里最好的初熟之物带到耶和华－你上帝的殿中。 “不可用母山羊的奶来煮它的小山羊。”
EXOD|23|20|“看哪，我要差遣使者在你前面，在路上保护你，领你到我所预备的地方。
EXOD|23|21|你们要在他面前谨慎，听从他的话。不可抗拒 他，否则他必不赦免你们的过犯，因为我的名在他身上。
EXOD|23|22|“你若真的听从他的话，照我一切所说的去做，我就以你的仇敌为仇敌，以你的敌人为敌人。
EXOD|23|23|“我的使者要走在你前面，领你到 亚摩利 人、 赫 人、 比利洗 人、 迦南 人、 希未 人、 耶布斯 人那里，我必将他们除灭。
EXOD|23|24|你不可跪拜事奉他们的神明，也不可随从他们的习俗，却要彻底废除，完全打碎他们的柱像。
EXOD|23|25|你们要事奉耶和华－你们的上帝，他必赐福给你的粮食和水，也必从你中间除去疾病。
EXOD|23|26|你境内必没有流产的、不生育的。我要使你享满你年日的数目。
EXOD|23|27|凡你所到的地方，我要使那里的众百姓在你面前惊慌失措，又要使你所有的仇敌转身逃跑。
EXOD|23|28|我要派瘟疫 在你的前面，把 希未 人、 迦南 人、 赫 人从你面前赶出去。
EXOD|23|29|我不在一年之内把他们从你面前赶出去，恐怕地会荒废，野地的走兽增多危害你。
EXOD|23|30|我要逐渐把他们从你面前赶出去，直到你的人数增多，承受那地为业。
EXOD|23|31|我要定你的疆界，从 红海 直到 非利士海 ，从旷野直到 大河 。我要把那地的居民交在你手中，你要把他们从你面前赶出去。
EXOD|23|32|不可跟他们和他们的神明立约。
EXOD|23|33|他们不可住在你的地上，免得他们使你得罪我。你若事奉他们的神明，必成为你的圈套。”
EXOD|24|1|耶和华对 摩西 说：“你和 亚伦 、 拿答 、 亚比户 ，以及 以色列 长老中的七十人，都要上到耶和华这里来，远远地下拜。
EXOD|24|2|只有 摩西 可以接近耶和华，其他的人却不可接近；百姓也不可和他一同上来。”
EXOD|24|3|摩西 下山，向百姓陈述耶和华一切的命令和典章。众百姓齐声说：“耶和华所吩咐的一切，我们都必遵行。”
EXOD|24|4|摩西 将耶和华一切的命令都写下来。 他清早起来，在山脚筑了一座坛，按着 以色列 十二支派立了十二根石柱。
EXOD|24|5|他差派 以色列 的年轻人去献燔祭，又宰牛献给耶和华为平安祭。
EXOD|24|6|摩西 将血的一半盛在盆中，另一半洒在坛上。
EXOD|24|7|然后，他拿起约书来，念给百姓听。他们说：“耶和华所吩咐的一切，我们都必遵行，也必听从。”
EXOD|24|8|摩西 把血洒在百姓身上，说：“看哪！这是立约的血，是耶和华按照这一切的命令和你们立约的凭据。”
EXOD|24|9|摩西 、 亚伦 、 拿答 、 亚比户 ，以及 以色列 长老中的七十人都上去，
EXOD|24|10|看见了 以色列 的上帝。在他的脚下，仿佛有蓝宝石铺道，明净如天。
EXOD|24|11|他不把手伸在 以色列 领袖的身上。他们瞻仰上帝，又吃又喝。
EXOD|24|12|耶和华对 摩西 说：“你上山到我这里来，就在那里，我要将石版，就是我所写的律法和诫命赐给你，使你可以教导他们。”
EXOD|24|13|摩西 和他的助手 约书亚 站起来； 摩西 上了上帝的山。
EXOD|24|14|摩西 对长老们说：“你们在这里等我们，直到我们再回到你们这里。看哪， 亚伦 和 户珥 与你们同在。谁有诉讼，可以去找他们。”
EXOD|24|15|摩西 上山，有云彩把山遮盖。
EXOD|24|16|耶和华的荣耀驻在 西奈山 ，云彩遮盖了山六天，第七天他从云中呼叫 摩西 。
EXOD|24|17|耶和华的荣耀在山顶上，在 以色列 人眼前，形状如吞噬的火。
EXOD|24|18|摩西 进入云中，登上了山。 摩西 在山上四十昼夜。
EXOD|25|1|耶和华吩咐 摩西 说：
EXOD|25|2|“你要吩咐 以色列 人献礼物给我。凡甘心乐意献给我的礼物，你们都可以收下。
EXOD|25|3|要从他们收的礼物是：金、银、铜，
EXOD|25|4|蓝色、紫色、朱红色纱 ，细麻，山羊毛，
EXOD|25|5|染红的公羊皮、精美的皮料，金合欢木，
EXOD|25|6|点灯的油，做膏油的香料、做香的香料，
EXOD|25|7|红玛瑙与宝石，可以镶嵌在以弗得和胸袋上。
EXOD|25|8|他们要为我造圣所，使我住在他们中间。
EXOD|25|9|你们要按照我指示你的，帐幕和其中一切器具的样式，照样去做。”
EXOD|25|10|“他们要用金合欢木做一个柜子，长二肘半，宽一肘半，高一肘半。
EXOD|25|11|你要把它里里外外包上纯金，四围要镶上金边。
EXOD|25|12|要铸造四个金环，安在柜子的四脚上；这边两个环，那边两个环。
EXOD|25|13|要用金合欢木做两根杠，包上金子。
EXOD|25|14|要把杠穿过柜旁的环，以便抬柜。
EXOD|25|15|这杠要留在柜的环内，不可抽出来。
EXOD|25|16|要把我所要赐给你的法版 放在柜里。
EXOD|25|17|要用纯金做一个柜盖 ，长二肘半，宽一肘半。
EXOD|25|18|要造两个用金子锤出的基路伯，从柜盖的两端锤出它们。
EXOD|25|19|这端锤出一个基路伯，那端锤出一个基路伯；从柜盖的两端锤出两个基路伯。
EXOD|25|20|二基路伯的翅膀要向上张开，用翅膀遮住柜盖，脸要彼此相对；基路伯的脸要朝向柜盖。
EXOD|25|21|要把柜盖安在柜的上边，又要把我所要赐给你的法版放在柜里。
EXOD|25|22|我要在那里与你相会，并要从法版之柜的柜盖上，两个基路伯的中间，将我要吩咐 以色列 人的一切事告诉你。”
EXOD|25|23|“你要用金合欢木做一张供桌，长二肘，宽一肘，高一肘半，
EXOD|25|24|把它包上纯金，四围镶上金边。
EXOD|25|25|供桌的四围各做一掌宽的边缘，边缘周围要镶上金边。
EXOD|25|26|要为供桌做四个金环，把环安在四个桌脚的四角上。
EXOD|25|27|环要靠近边缘，以便穿杠抬供桌。
EXOD|25|28|要用金合欢木做两根杠，包上金子，用来抬供桌。
EXOD|25|29|要用纯金做桌上的盘、碟，以及浇酒祭的壶和杯。
EXOD|25|30|要把供饼摆在桌上，常在我面前。”
EXOD|25|31|“要造一座用纯金锤出的灯台。灯台的座、干、杯、花萼和花瓣，都要和灯台接连一块。
EXOD|25|32|灯台两旁要伸出六根枝子：这边三根，那边三根。
EXOD|25|33|这边枝子上有三个杯，形状像杏花，有花萼有花瓣；那边枝子上也有三个杯，形状像杏花，有花萼有花瓣。从灯台伸出来的六根枝子都是如此。
EXOD|25|34|灯台本身要有四个杯，形状像杏花，有花萼有花瓣。
EXOD|25|35|灯台的第一对枝子下面有花萼，灯台的第二对枝子下面有花萼，灯台的第三对枝子下面也有花萼；灯台伸出的六根枝子都是如此。
EXOD|25|36|花萼和枝子都要和灯台接连一块，全是从一块纯金锤出来的。
EXOD|25|37|要做灯台的七盏灯，灯要点燃，照亮前面。
EXOD|25|38|要用纯金做灯剪和灯盘。
EXOD|25|39|做灯台和这一切的器具要用一他连得纯金。
EXOD|25|40|要谨慎，照着在山上指示你的样式去做。”
EXOD|26|1|“你要用十幅幔子做帐幕。这些幔子要用搓的细麻和蓝色、紫色、朱红色纱织成，并且以刺绣的手艺绣上基路伯。
EXOD|26|2|每幅幔子要长二十八肘，每幅幔子宽四肘，全部的幔子尺寸都要一样。
EXOD|26|3|这五幅幔子要彼此相连；那五幅也彼此相连。
EXOD|26|4|在这一组相连幔子的末幅边上要缝蓝色的钮环；在另一组相连幔子的末幅边上也要照样做。
EXOD|26|5|这幅幔子上要缝五十个钮环，另一组相连幔子的末幅上也缝五十个钮环，环环相对。
EXOD|26|6|要做五十个金钩，用钩子使幔子彼此相连，成为一个帐幕。
EXOD|26|7|“你要用山羊毛织十一幅幔子来作帐幕的罩棚。
EXOD|26|8|每幅幔子要长三十肘，每幅幔子宽四肘；十一幅幔子的尺寸都要一样。
EXOD|26|9|要把五幅幔子连成一幅，又把六幅幔子连成一幅，这第六幅幔子要在罩棚的前面摺上去。
EXOD|26|10|在这一组相连幔子的末幅边上要缝五十个钮环；在另一组相连幔子的末幅边上也缝五十个钮环。
EXOD|26|11|要做五十个铜钩，钩在钮环中，使罩棚相连成为一个。
EXOD|26|12|罩棚幔子余下垂着的，那余下的半幅要垂在帐幕的背面。
EXOD|26|13|罩棚的幔子两旁所余下的，这边一肘，那边一肘，要垂在帐幕的两边，盖住帐幕。
EXOD|26|14|要用染红的公羊皮做罩棚的盖，再用精美皮料做外层的盖。
EXOD|26|15|“你要用金合欢木做竖立帐幕的木板，
EXOD|26|16|木板要长十肘，每块板宽一肘半，
EXOD|26|17|每块板有两个榫头可以彼此衔接。帐幕一切的板都要这样做。
EXOD|26|18|你要做帐幕的木板：南面，就是面向南方的那一边，要做二十块板。
EXOD|26|19|在这二十块板底下要做四十个带卯眼的银座；两个卯眼接连这块板上的两个榫头，另外两个卯眼接连那块板上的两个榫头。
EXOD|26|20|帐幕的第二边，就是北面，也要做二十块板，
EXOD|26|21|和四十个带卯眼的银座；这块板底下有两个卯眼，那块板底下也有两个卯眼。
EXOD|26|22|帐幕的后面，就是西面，要做六块板。
EXOD|26|23|帐幕后面的角落要做两块板。
EXOD|26|24|下端的板是成双的，上端要连在一起，直到顶端的第一个环子；两块板都要这样，做成两个角落。
EXOD|26|25|一共有八块板和十六个带卯眼的银座；这块板底下有两个卯眼，那块板底下也有两个卯眼。
EXOD|26|26|“你要用金合欢木做横木：为帐幕这面的板做五根横木，
EXOD|26|27|为帐幕那面的板做五根横木，又为帐幕后面，就是朝西的板做五根横木。
EXOD|26|28|板腰间的横木，要从一头通到另一头。
EXOD|26|29|板要包上金子，又要做板上的金环来套横木；横木也要包上金子。
EXOD|26|30|要照着在山上所指示你的样式，把帐幕竖立起来。
EXOD|26|31|“你要用蓝色、紫色、朱红色纱，和搓的细麻织幔子，以刺绣的手艺绣上基路伯。
EXOD|26|32|要把幔子挂在四根包金的金合欢木柱子上，柱子有金钩，并且安在四个带卯眼的银座上。
EXOD|26|33|要把幔子垂挂在钩子上，把法柜抬进幔子内；这幔子要将圣所和至圣所隔开。
EXOD|26|34|又要把柜盖安在至圣所内的法柜上，
EXOD|26|35|把供桌安在幔子的外面，供桌在北面，灯台在帐幕的南面，和供桌相对。
EXOD|26|36|“你要用蓝色、紫色、朱红色纱，和搓的细麻，以刺绣的手艺为帐幕织门帘。
EXOD|26|37|要用金合欢木为帘子做五根柱子，包上金子。柱子有金钩，又为柱子铸造五个带卯眼的铜座。”
EXOD|27|1|“你要用金合欢木做祭坛，长五肘，宽五肘，这坛是正方形的，高三肘。
EXOD|27|2|要在坛的四角做四个翘角，与坛接连一块；要把坛包上铜。
EXOD|27|3|要做桶子来盛坛上的灰，又要做铲子、盘子、肉叉和火盆；坛上一切的器具都要用铜做。
EXOD|27|4|要为坛做一个铜网，在网的四角做四个铜环，
EXOD|27|5|把网安在坛四围的边的下面，使网垂到坛的半腰。
EXOD|27|6|又要用金合欢木为坛做杠，包上铜。
EXOD|27|7|这杠要穿过坛两旁的环子，用来抬坛。
EXOD|27|8|要用板做坛，坛的中心是空的，都照着在山上所指示你的样式做。”
EXOD|27|9|“你要做帐幕的院子。南面，就是面向南方的那一边，要用搓的细麻做院子的帷幔，长一百肘，
EXOD|27|10|院子要有二十根柱子，二十个带卯眼的铜座。要用银做柱子的钩和箍。
EXOD|27|11|北面的长度也一样，帷幔长一百肘，要有二十根柱子，二十个带卯眼的铜座。要用银做柱子的钩和箍。
EXOD|27|12|院子的西面有帷幔，宽五十肘，帷幔要有十根柱子，十个带卯眼的座。
EXOD|27|13|院子的东面，就是面向东方的那一边，宽五十肘。
EXOD|27|14|一边的帷幔有十五肘，要有三根柱子，三个带卯眼的座。
EXOD|27|15|另一边的帷幔也有十五肘，要有三根柱子，三个带卯眼的座。
EXOD|27|16|院子的门要有二十肘长的帘子，用蓝色、紫色、朱红色纱，和搓的细麻，以刺绣的手艺织成；要有四根柱子，四个带卯眼的座。
EXOD|27|17|院子四围一切的柱子都要用银子箍着，要用银做柱子的钩子，用铜做带卯眼的座。
EXOD|27|18|院子要长一百肘，宽五十肘 ，高五肘。要用搓的细麻做帷幔，用铜做带卯眼的座。
EXOD|27|19|帐幕中各样用途的器具，以及帐幕一切的橛子和院子里一切的橛子，都要用铜做。”
EXOD|27|20|“你要吩咐 以色列 人，把捣成的纯橄榄油拿来给你，用以点灯，使灯经常点着；
EXOD|27|21|在会幕中法柜前的幔子外， 亚伦 和他的儿子要从晚上到早晨，在耶和华面前照管这灯。这要成为 以色列 人世世代代永远的定例。”
EXOD|28|1|“你要从 以色列 人中，叫你的哥哥 亚伦 和他的儿子 拿答 、 亚比户 、 以利亚撒 、 以他玛 一同亲近你，作事奉我的祭司。
EXOD|28|2|你要为你哥哥 亚伦 做圣衣，以示尊严和华美。
EXOD|28|3|要吩咐一切心中有智慧的，就是我用智慧的灵所充满的人，为 亚伦 做衣服，使他分别为圣，作事奉我的祭司。
EXOD|28|4|所要做的是胸袋、以弗得、外袍、织成的内袍、礼冠和腰带。他们要为你哥哥 亚伦 和他的儿子做圣衣，使他们作祭司事奉我。
EXOD|28|5|要用金色、蓝色、紫色、朱红色纱，和细麻去缝制。
EXOD|28|6|“他们要用金色、蓝色、紫色、朱红色纱，和搓的细麻，以刺绣的手艺做以弗得。
EXOD|28|7|以弗得当有两条肩带，接上两端，使它相连。
EXOD|28|8|以弗得的精致带子，要以一样的手艺，用金色、蓝色、紫色、朱红色纱，和搓的细麻缝制，与以弗得接连在一起。
EXOD|28|9|要取两块红玛瑙，在上面刻 以色列 儿子的名字：
EXOD|28|10|六个名字在一块宝石上，六个名字在另一块宝石上，都按照他们出生的次序。
EXOD|28|11|要以雕刻宝石的手艺，如同刻印章，把 以色列 儿子的名字刻在这两块宝石上，并把宝石镶在金槽里。
EXOD|28|12|要把这两块宝石安在以弗得的两条肩带上，为 以色列 人作纪念石。 亚伦 要在耶和华面前把他们的名字带在两肩上，作为纪念。
EXOD|28|13|要用金子做两个槽，
EXOD|28|14|再用纯金打两条链子，像编成的绳子一样，把这编成的金链扣在槽上。”
EXOD|28|15|“你要以刺绣的手艺做一个决断的胸袋，和做以弗得的方法一样，用金色、蓝色、紫色、朱红色纱，和搓的细麻缝制。
EXOD|28|16|胸袋是正方形的，叠成两层，长一虎口，宽一虎口。
EXOD|28|17|要在上面镶四行宝石：第一行是红宝石、红璧玺、红玉；
EXOD|28|18|第二行是绿宝石、蓝宝石、金刚石；
EXOD|28|19|第三行是紫玛瑙、白玛瑙、紫晶；
EXOD|28|20|第四行是水苍玉、红玛瑙、碧玉。这些都要镶在金槽中。
EXOD|28|21|这些宝石要有 以色列 十二个儿子的名字，如同刻印章，每一颗有自己的名字，代表十二个支派。
EXOD|28|22|要在胸袋上用纯金打链子，像编成的绳子一样。
EXOD|28|23|要为胸袋做两个金环，把这两个环安在胸袋的两端。
EXOD|28|24|要把那两条编成的金链系在胸袋两端的两个环上。
EXOD|28|25|又要把链子的另外两端扣在两个槽上，安在以弗得前面的肩带上。
EXOD|28|26|要做两个金环，安在胸袋的两端，在以弗得里面的边上。
EXOD|28|27|再做两个金环，安在以弗得前面两条肩带的下边，靠近接缝处，在以弗得精致带子的上面。
EXOD|28|28|要用蓝色的带子把胸袋的环与以弗得的环系住，使胸袋绑在以弗得的精致带子上，不致松脱。
EXOD|28|29|亚伦 进圣所的时候，要把刻着 以色列 儿子名字的决断胸袋带着，放在心上，在耶和华面前常作纪念。
EXOD|28|30|又要将乌陵和土明 放在决断胸袋里； 亚伦 进到耶和华面前的时候，要放在心上。这样， 亚伦 在耶和华面前要把 以色列 人的决断胸袋常常带着，放在心上。”
EXOD|28|31|“你要做以弗得的外袍，颜色全是蓝的。
EXOD|28|32|袍上方的中间要留一个领口，领口周围的领边要以手艺编织而成，好像铠甲的领口，免得破裂。
EXOD|28|33|袍子下摆，就是下摆的周围要用蓝色、紫色、朱红色纱做石榴，周围的石榴中间要有金铃铛：
EXOD|28|34|一个金铃铛一个石榴，一个金铃铛一个石榴，在袍子下摆的周围。
EXOD|28|35|亚伦 供职的时候要穿这袍。他进入圣所到耶和华面前，以及出来的时候，袍上的铃声必被听见，使他不至于死。
EXOD|28|36|“你要用纯金做一面牌，如同刻印章，在上面刻‘归耶和华为圣’。
EXOD|28|37|要用蓝色的带子把牌系在礼冠上，在礼冠的正前面。
EXOD|28|38|这牌必在 亚伦 的额上， 亚伦 要担当干犯圣物的罪孽；这圣物是 以色列 人在一切圣礼物上所分别为圣的。这牌要常在他的额上，使他们可以在耶和华面前蒙悦纳。
EXOD|28|39|要用细麻编织内袍，用细麻做礼冠，又以刺绣的手艺做腰带。
EXOD|28|40|“你要为 亚伦 的儿子做内袍、腰带、头巾，以示尊严和华美。
EXOD|28|41|要把这些给你哥哥 亚伦 和他的儿子穿戴，又要膏他们，授予圣职，使他们分别为圣，作事奉我的祭司。
EXOD|28|42|要用细麻布给他们做裤子来遮掩下体，从腰间直到大腿。
EXOD|28|43|亚伦 和他儿子进入会幕，或接近祭坛，在圣所供职的时候要穿上裤子，免得担当罪孽而死。这要成为 亚伦 和他后裔永远的定例。”
EXOD|29|1|“这是你使他们分别为圣，作事奉我的祭司时要做的事：取一头公牛犊，两只无残疾的公绵羊，
EXOD|29|2|无酵饼、用油调和的无酵饼，和抹油的无酵薄饼；这些饼都要用细麦面做成。
EXOD|29|3|这些饼要装在一个篮子里，用篮子带来，又把公牛和两只公绵羊牵来。
EXOD|29|4|要带 亚伦 和他儿子到会幕的门口，用水洗他们。
EXOD|29|5|要拿服装，给 亚伦 穿上内袍和以弗得的外袍，以及以弗得，又带上胸袋，束上以弗得精致的带子。
EXOD|29|6|要把礼冠戴在他头上，将圣冕加在礼冠上，
EXOD|29|7|把膏油倒在他头上膏他。
EXOD|29|8|要带他的儿子来，给他们穿上内袍。
EXOD|29|9|要给 亚伦 和他的儿子束上腰带，裹上头巾，他们就凭永远的定例得祭司的职分。又要授圣职给 亚伦 和他的儿子。
EXOD|29|10|“你要把公牛牵到会幕前， 亚伦 和他的儿子要按手在公牛的头上。
EXOD|29|11|你要在耶和华面前，在会幕的门口宰这公牛。
EXOD|29|12|要取些公牛的血，用指头抹在祭坛的四个翘角上，把其余的血全倒在坛的底座上。
EXOD|29|13|要把所有包着内脏的脂肪、肝上的网油、两个肾和肾上的脂肪，都烧在坛上。
EXOD|29|14|只是公牛的肉、皮、粪都要在营外用火焚烧；这牛是赎罪祭。
EXOD|29|15|“你要牵一只公绵羊来， 亚伦 和他儿子要按手在这羊的头上。
EXOD|29|16|你要宰这羊，把血洒在祭坛的周围。
EXOD|29|17|再把羊切成肉块，洗净内脏和腿，连肉块和头放在一处。
EXOD|29|18|要把全羊烧在坛上。这是献给耶和华的燔祭，是献给耶和华馨香的火祭。”
EXOD|29|19|“你要把第二只公绵羊牵来， 亚伦 和他儿子要按手在这羊的头上。
EXOD|29|20|你要宰这羊，取些血抹在 亚伦 的右耳垂和他儿子的右耳垂上，又抹在他们右手的大拇指和右脚的大脚趾上，然后把其余的血洒在坛的周围。
EXOD|29|21|你要取些膏油和坛上的血，弹在 亚伦 和他的衣服上，以及他儿子和他们的衣服上； 亚伦 和他的衣服，他儿子和他们的衣服都成为圣了。
EXOD|29|22|“你要取这羊的脂肪，肥尾巴、包着内脏的脂肪、肝上的网油、两个肾、肾上的脂肪和右腿，这是圣职礼所献的公绵羊；
EXOD|29|23|再从耶和华面前那装无酵饼的篮子中取一个饼、一个油饼和一个薄饼，
EXOD|29|24|把它们都放在 亚伦 的手和他儿子的手上，在耶和华面前摇一摇，作为摇祭。
EXOD|29|25|然后，你要从他们手中接过来，放在燔祭上，一起烧在坛上，作为耶和华面前馨香之气；这是献给耶和华的火祭。
EXOD|29|26|“你要取 亚伦 圣职礼所献公绵羊的胸，在耶和华面前摇一摇，作为摇祭；这份就是你的。
EXOD|29|27|那摇祭的胸和举祭的腿，就是圣职礼献公绵羊时所摇的、所举的，你要使它们分别为圣，是归给 亚伦 和他儿子的。
EXOD|29|28|这是 亚伦 和他子孙凭永远的定例从 以色列 人中所应得的；因为这是举祭，是从 以色列 人的平安祭中取出，作为献给耶和华的举祭。
EXOD|29|29|“ 亚伦 的圣衣要传给他的子孙，使他们在受膏和承接圣职的时候穿上。
EXOD|29|30|他的子孙接续他当祭司的，每逢进入会幕在圣所供职的时候，要穿这圣衣七天。
EXOD|29|31|“你要拿圣职礼所献的公绵羊，在圣处煮它的肉。
EXOD|29|32|亚伦 和他儿子要在会幕的门口吃这羊的肉和篮子里的饼。
EXOD|29|33|他们要吃那些用来赎罪之物，好承接圣职，使他们分别为圣。外人不可吃，因为这是圣物。
EXOD|29|34|那圣职礼所献的肉或饼，若有剩余留到早晨，就要把剩下的用火烧了，不可再吃，因为这是圣物。
EXOD|29|35|“你要这样照我一切所吩咐的，向 亚伦 和他儿子行授圣职礼七天。
EXOD|29|36|为了赎罪，每天要献一头公牛为赎罪祭。你要为祭坛赎罪，使坛洁净，并要用膏抹坛，使坛成为圣。
EXOD|29|37|要为坛赎罪七天，使坛成为圣，坛就成为至圣。凡触摸坛的都成为圣。”
EXOD|29|38|“这是你要献在坛上的：每天不可间断地献两只一岁的羔羊；
EXOD|29|39|早晨献第一只羔羊，黄昏献第二只羔羊。
EXOD|29|40|献第一只羔羊时，要同时献上十分之一伊法细面，调和四分之一欣捣成的油，再献四分之一欣酒作浇酒祭。
EXOD|29|41|黄昏你献第二只羔羊，要照早晨的素祭和同献的浇酒祭献上，作为献给耶和华馨香的火祭。
EXOD|29|42|这要在耶和华面前，在会幕的门口，作为你们世世代代经常献的燔祭。我要在那里与你们 相会，和你说话。
EXOD|29|43|我要在那里与 以色列 人相会，会幕就要因我的荣耀成为圣。
EXOD|29|44|我要使会幕和祭坛分别为圣，也要使 亚伦 和他的儿子分别为圣，作事奉我的祭司。
EXOD|29|45|我要住在 以色列 人中，作他们的上帝。
EXOD|29|46|他们必知道我是耶和华－他们的上帝，是将他们从 埃及 地领出来的，为要住在他们中间。我是耶和华－他们的上帝 。”
EXOD|30|1|“你要用金合欢木做一座烧香的坛，
EXOD|30|2|长一肘，宽一肘，这坛是正方形的，高二肘。坛的四个翘角与坛接连一块。
EXOD|30|3|要把坛的上面与坛的四围，以及坛的四个翘角包上纯金；又要在坛的四围镶上金边。
EXOD|30|4|要在坛的两个对侧，金边下面做两个金环，用来穿杠抬坛。
EXOD|30|5|要用金合欢木做杠，包上金子。
EXOD|30|6|要把坛放在法柜前的幔子外，对着法柜上的柜盖，就是我与你相会的地方。
EXOD|30|7|亚伦 要在坛上烧芬芳的香；每早晨整理灯的时候，他都要烧这香。
EXOD|30|8|黄昏点灯的时候， 亚伦 也要烧这香。这是你们世世代代在耶和华面前常烧的香。
EXOD|30|9|在这坛上不可烧别样的香，不可献燔祭、素祭，也不可献浇酒祭。
EXOD|30|10|亚伦 每年一次要为坛的四个翘角赎罪。他每年一次要用赎罪祭的血为坛赎罪，作为世世代代的定例。这坛在耶和华面前是至圣的。”
EXOD|30|11|耶和华吩咐 摩西 说：
EXOD|30|12|“你数点 以色列 人，计算人头时，被数的每一个人要把他生命的赎价献给耶和华，免得灾殃在数点中临到他们。
EXOD|30|13|每一个被数的人要按照圣所的舍客勒，付半舍客勒，一舍客勒是二十季拉；这半舍客勒是献给耶和华的礼物。
EXOD|30|14|每一个被数的人，就是二十岁以上的，要将这礼物献给耶和华。
EXOD|30|15|富有的不必多付，贫穷的也不可少出，各人都要献半舍客勒给耶和华，作你们生命的赎价。
EXOD|30|16|你要向 以色列 人收这赎罪的银子，用在会幕的事工。这要在耶和华面前为 以色列 人作纪念，作你们生命的赎价。”
EXOD|30|17|耶和华吩咐 摩西 说：
EXOD|30|18|“你要用铜做洗濯盆和盆座，用来洗濯。要将盆放在会幕和祭坛的中间，盆里盛水。
EXOD|30|19|亚伦 和他的儿子要用这盆洗手洗脚。
EXOD|30|20|他们进会幕，或是走近坛前供职，献火祭给耶和华的时候，必须用水洗濯，免得死亡；
EXOD|30|21|他们要洗手洗脚，免得死亡。这是 亚伦 和他的后裔世世代代永远的定例。”
EXOD|30|22|耶和华吩咐 摩西 说：
EXOD|30|23|“你要取上等的香料，就是五百舍客勒流质的没药、二百五十香肉桂、二百五十香菖蒲，
EXOD|30|24|和五百桂皮，都按照圣所的舍客勒；再取一欣橄榄油，
EXOD|30|25|以做香的方法调和制成圣膏油，它就成为圣膏油。
EXOD|30|26|要用这膏油抹会幕和法柜，
EXOD|30|27|供桌和供桌的一切器具，灯台和灯台的器具 ，以及香坛、
EXOD|30|28|燔祭坛和坛的一切器具，洗濯盆和盆座。
EXOD|30|29|你要使这些分别为圣，成为至圣；凡触摸它们的都成为圣。
EXOD|30|30|要膏 亚伦 和他的儿子，使他们分别为圣，作事奉我的祭司。
EXOD|30|31|你要吩咐 以色列 人说：‘你们要世世代代以这油为我的圣膏油。
EXOD|30|32|不可把这油倒在别人身上，也不可用配制这膏油的方法制成同样的膏油。这膏油是圣的，你们要以它为圣。
EXOD|30|33|凡调和与此类似的膏油，或将它膏在别人身上的，这人要从百姓中剪除。’”
EXOD|30|34|耶和华吩咐 摩西 说：“你要取香料，就是拿他弗、施喜列、喜利比拿，这些香料再加纯乳香，每样都要相同的分量。
EXOD|30|35|你要用这些加上盐，以配制香料的方法，制成纯净又神圣的香。
EXOD|30|36|要取一点这香，捣成细的粉，放在会幕中的法柜前，就是我和你相会的地方。你们要以这香为至圣。
EXOD|30|37|你们不可用这配制的方法为自己做香；要以这香为圣，归于耶和华。
EXOD|30|38|为要闻香味而配制同样的香的，这人要从百姓中剪除。”
EXOD|31|1|耶和华吩咐 摩西 说：
EXOD|31|2|“你看，我已经题名召 犹大 支派中 户珥 的孙子， 乌利 的儿子 比撒列 。
EXOD|31|3|我以上帝的灵充满他，使他有智慧，有聪明，有知识，能做各样的工，
EXOD|31|4|能设计图案，用金、银、铜制造各物，
EXOD|31|5|又能雕刻镶嵌用的宝石，雕刻木头，做各样的工。
EXOD|31|6|看哪，我委派 但 支派中 亚希撒抹 的儿子 亚何利亚伯 与他同工。凡心里有智慧的，我更要赐给他们智慧的心，能做我所吩咐你的一切，
EXOD|31|7|就是会幕、法柜和其上的柜盖、会幕中一切的器具、
EXOD|31|8|供桌和供桌的器具、纯金的灯台和灯台的一切器具、香坛、
EXOD|31|9|燔祭坛和坛的一切器具、洗濯盆与盆座、
EXOD|31|10|供祭司职分用的精致礼服， 亚伦 祭司的圣衣和他儿子的衣服，
EXOD|31|11|以及膏油和圣所用的芬芳的香。他们都要照我所吩咐的一切去做。”
EXOD|31|12|耶和华对 摩西 说：
EXOD|31|13|“你要吩咐 以色列 人说：‘你们务要守我的安息日，因为这是你我之间世世代代的记号，叫你们知道我是耶和华，是使你们分别为圣的。
EXOD|31|14|你们要守安息日，以它为圣日。凡干犯这日的，必被处死；凡在这日做工的，那人必从百姓中剪除。
EXOD|31|15|六日要做工，但第七日是向耶和华守完全安息的安息圣日。凡在安息日做工的，必被处死。’
EXOD|31|16|以色列 人要守安息日，世世代代守安息日为永远的约。
EXOD|31|17|这是我和 以色列 人之间永远的记号，因为六日之内耶和华造天地，第七日就安息舒畅。”
EXOD|31|18|耶和华在 西奈山 和 摩西 说完了话，就把两块法版交给他，是上帝用指头写的石版。
EXOD|32|1|百姓见 摩西 迟迟不下山，就聚集到 亚伦 那里，对他说：“起来！为我们造神明，在我们前面引路，因为领我们出 埃及 地的那个 摩西 ，我们不知道他遭遇了什么事。”
EXOD|32|2|亚伦 对他们说：“你们去摘下你们妻子、儿女耳上的金环，拿来给我。”
EXOD|32|3|众百姓就摘下他们耳上的金环，拿来给 亚伦 。
EXOD|32|4|亚伦 从他们手里接过来，用模子塑造它，把它铸成一头牛犊。他们就说：“ 以色列 啊，这是领你出 埃及 地的神明！”
EXOD|32|5|亚伦 看见，就在牛犊面前筑坛。 亚伦 宣告说：“明日要向耶和华守节。”
EXOD|32|6|次日清早，百姓起来献燔祭和平安祭，就坐下吃喝，起来玩乐。
EXOD|32|7|耶和华吩咐 摩西 ：“下去吧，因为你从 埃及 领上来的百姓已经败坏了。
EXOD|32|8|他们这么快偏离了我所吩咐的道，为自己铸了一头牛犊，向它跪拜，向它献祭，说：‘ 以色列 啊，这就是领你出 埃及 地的神明。’”
EXOD|32|9|耶和华对 摩西 说：“我看这百姓，看哪，他们真是硬着颈项的百姓。
EXOD|32|10|现在，你且由着我，我要向他们发烈怒，灭绝他们，但我要使你成为大国。”
EXOD|32|11|摩西 就恳求耶和华－他的上帝，说：“耶和华啊，你为什么向你的百姓发烈怒呢？这百姓是你用大能大力的手从 埃及 地领出来的！
EXOD|32|12|为什么让 埃及 人说：‘他领他们出去，是要降灾祸给他们，在山中把他们杀了，将他们从地上除灭’呢？求你回心转意，不发你的烈怒，不降灾祸给你的百姓。
EXOD|32|13|求你记念你的仆人 亚伯拉罕 、 以撒 、 以色列 。你曾向他们指着自己起誓说：‘我必使你们的后裔像天上的星那样多，并且我要将所应许的这全地赐给你们的后裔，让他们永远承受为业。’”
EXOD|32|14|于是耶和华改变心意，不把所说的灾祸降给他的百姓。
EXOD|32|15|摩西 转身下山，手里拿着两块法版。这版的两面都写着字，正面背面都有字。
EXOD|32|16|版是上帝的工作，字是上帝写的字，刻在版上。
EXOD|32|17|约书亚 一听见百姓呼喊的声音，就对 摩西 说：“在营里有战争的声音。”
EXOD|32|18|摩西 说：“这不是打胜仗的声音，也不是打败仗的声音，我听见的是歌唱的声音。”
EXOD|32|19|摩西 走近营前，看见牛犊，又看见人在跳舞，就发烈怒，把两块版从手中扔到山下摔碎了。
EXOD|32|20|他将他们所铸的牛犊用火焚烧，磨得粉碎，撒在水面上，叫 以色列 人喝。
EXOD|32|21|摩西 对 亚伦 说：“这百姓向你做了什么呢？你竟使他们陷入大罪中！”
EXOD|32|22|亚伦 说：“求我主不要发烈怒。你知道这百姓，他们是向恶的。
EXOD|32|23|他们对我说：‘你为我们造神明，在我们前面引路，因为领我们出 埃及 地的那个 摩西 ，我们不知道他遭遇了什么事。’
EXOD|32|24|我对他们说：‘凡有金环的可以摘下来’，他们就给了我。我把金环扔在火中，这牛犊就出来了。”
EXOD|32|25|摩西 见百姓放肆，因 亚伦 纵容他们，使这事成了敌人的笑柄，
EXOD|32|26|就站在营门前，说：“凡属耶和华的人，都到我这里来！”于是 利未 人都聚集到他那里。
EXOD|32|27|他对他们说：“耶和华－ 以色列 的上帝这样说：‘你们各人把刀佩在腰间，从这门到那门，来回走遍全营，各人要杀自己的弟兄、邻舍和亲人。’”
EXOD|32|28|利未 人遵照 摩西 的话做了。那一天百姓中倒下的约有三千人。
EXOD|32|29|摩西 说：“今天你们要奉献自己 来事奉耶和华，因为各人牺牲自己的儿子和弟兄，使耶和华今天赐福给你们。”
EXOD|32|30|第二天， 摩西 对百姓说：“你们犯了大罪。我如今要上耶和华那里去，或许可以为你们赎罪。”
EXOD|32|31|摩西 回到耶和华那里，说：“唉！这百姓犯了大罪，为自己造了金的神明。
EXOD|32|32|现在，求你赦免他们的罪；不然，就把我从你所写的册上除名。”
EXOD|32|33|耶和华对 摩西 说：“谁得罪我，我就把他从我的册上除去。
EXOD|32|34|现在你去，领这百姓往我所告诉你的地方去，看哪，我的使者必在你的前面引路。到了该惩罚的时候，我必惩罚他们的罪。”
EXOD|32|35|耶和华降灾与百姓，因为他们和 亚伦 一起造了牛犊。
EXOD|33|1|耶和华吩咐 摩西 说：“去，离开这里，你和你从 埃及 地领出来的百姓要上到我起誓应许给 亚伯拉罕 、 以撒 和 雅各 之地去；我曾对他们说：‘我要将这地赐给你的后裔’。
EXOD|33|2|我要差遣使者在你前面，把 迦南 人、 亚摩利 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人赶出
EXOD|33|3|那流奶与蜜之地。但我不与你们上去，因为你们是硬着颈项的百姓，免得我在路上把你们灭绝。”
EXOD|33|4|百姓一听见这坏的信息，他们就悲哀，没有人佩戴首饰。
EXOD|33|5|耶和华对 摩西 说：“你对 以色列 人说：‘你们是硬着颈项的百姓，我若在你们中间一起上去，只一瞬间，就必把你们灭绝。现在把你们身上的首饰摘下来，我好知道该怎样处置你们。’”
EXOD|33|6|以色列 人离开 何烈山 以后，就把身上的首饰全都摘下来。
EXOD|33|7|摩西 拿一个帐棚支搭在营外，离营有一段距离，他称这帐棚为会幕。凡求问耶和华的，就到营外的会幕那里去。
EXOD|33|8|当 摩西 出营到会幕去的时候，百姓就都起来，各人站在自己帐棚的门口，望着 摩西 ，直到他进了会幕。
EXOD|33|9|摩西 进会幕的时候，云柱就降下来，停在会幕的门前，耶和华就与 摩西 说话。
EXOD|33|10|众百姓看见云柱停在会幕的门前，就都起来，各人在自己帐棚的门口下拜。
EXOD|33|11|耶和华与 摩西 面对面说话，好像人与朋友说话。 摩西 回到营里去，他的年轻助手 嫩 的儿子 约书亚 却没有离开会幕。
EXOD|33|12|摩西 对耶和华说：“看，你曾对我说：‘将这百姓领上去’；却没有让我知道你要差派谁与我同去。你还说：‘我按你的名认识你，你也在我眼前蒙了恩。’
EXOD|33|13|我如今若在你眼前蒙恩，求你将你的道指示我，使我可以认识你，并在你眼前蒙恩。求你顾念这国是你的子民。”
EXOD|33|14|耶和华说：“我必亲自去，让你安心。”
EXOD|33|15|摩西 说：“你若不亲自去，就不要把我们从这里领上去。
EXOD|33|16|现在，人如何得知我和你的百姓在你眼前蒙恩呢？岂不是因为你与我们同去，使我和你的百姓与地面上的万民有分别吗？”
EXOD|33|17|耶和华对 摩西 说：“你所说的这件事，我也会去做，因为你在我眼前蒙了恩，并且我按你的名认识你。”
EXOD|33|18|摩西 说：“求你显出你的荣耀给我看。”
EXOD|33|19|耶和华说：“我要显示我一切的美善，在你面前经过，并要在你面前宣告耶和华的名。我要恩待谁就恩待谁，要怜悯谁就怜悯谁。”
EXOD|33|20|他又说：“只是你不能看见我的面，因为没有人看见我还可以存活。”
EXOD|33|21|耶和华说：“看哪，靠近我这里有个地方，你可以站在这磐石上。
EXOD|33|22|当我的荣耀经过的时候，我必将你放在磐石缝里，用我的手掌遮掩你，等我过去，
EXOD|33|23|然后我要将我的手掌收回，你就可以看见我的背，却看不到我的面。”
EXOD|34|1|耶和华对 摩西 说：“你要凿出两块石版，和先前的一样；我要把你摔碎的那版上先前所写的字，写在这版上。
EXOD|34|2|明日早晨，你要预备好了，上 西奈山 ，在山顶那里站在我面前。
EXOD|34|3|谁也不可和你上去，整座山都不可见到人，也不可有羊群牛群在山下吃草。”
EXOD|34|4|摩西 就凿出两块石版，和先前的一样。他清晨起来，遵照耶和华吩咐他的，上 西奈山 去，手里拿着两块石版。
EXOD|34|5|耶和华在云中降临，与 摩西 一同站在那里，宣告耶和华的名。
EXOD|34|6|耶和华在他面前经过，宣告： “耶和华，耶和华， 有怜悯，有恩惠的上帝， 不轻易发怒， 且有丰盛的慈爱和信实，
EXOD|34|7|为千代的人存留慈爱， 赦免罪孽、过犯和罪恶， 万不以有罪的为无罪， 必惩罚人的罪， 自父及子，直到三、四代。”
EXOD|34|8|摩西 急忙俯伏在地敬拜，
EXOD|34|9|说：“主啊，我若在你眼前蒙恩，求主在我们中间同行。虽然这是硬着颈项的百姓，求你赦免我们的罪孽和罪恶，接纳我们为你的产业。”
EXOD|34|10|耶和华说：“看哪，我要立约，要在你众百姓面前行奇妙的事，是在全地万国中未曾做过的。你周围的万民要看见我藉着你所行，耶和华可畏惧的作为。
EXOD|34|11|“我今天所吩咐你的，你要谨守。看哪，我要从你面前赶出 亚摩利 人、 迦南 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人。
EXOD|34|12|你要谨慎，不可与你所要去那地的居民立约，免得他们成为你中间的圈套。
EXOD|34|13|你要拆毁他们的祭坛，打碎他们的柱像，砍断他们的 亚舍拉 。
EXOD|34|14|不可敬拜别神，因为耶和华是忌邪 的上帝，他的名是忌邪者。
EXOD|34|15|你不可与那地的居民立约，因为他们随从自己的神明行淫；祭他们神明的时候，有人邀请你参加，你就会吃他的祭物。
EXOD|34|16|你为你儿子娶他们的女儿为妻，他们的女儿因着随从她们的神明行淫，就引诱你的儿子也随从她们的神明行淫。
EXOD|34|17|“不可为自己铸造神像。
EXOD|34|18|“你要守除酵节，照我所吩咐你的，在亚笔月内所定的日期吃无酵饼七天，因为你是在亚笔月内出了 埃及 。
EXOD|34|19|“凡头生的都是我的；无论是牛是羊，一切头生的公的牲畜都要分别出来 。
EXOD|34|20|头生的驴可以用羔羊代赎。若不赎它，就要打断它的颈项。凡头生的儿子都要赎出来。没有人可以空手来朝见我。
EXOD|34|21|“六日你要做工，第七日要安息，即使在耕种或收割的时候也要安息。
EXOD|34|22|在收割初熟麦子的时候要守七七节，又要在年底守收藏节。
EXOD|34|23|你所有的男丁要一年三次朝见主耶和华－ 以色列 的上帝。
EXOD|34|24|我要从你面前赶走列国，扩张你的疆界。你一年三次上去朝见耶和华－你上帝的时候，必没有人贪图你的地。
EXOD|34|25|“不可将我祭牲的血和有酵之物一同献上。逾越节的祭牲也不可留到早晨。
EXOD|34|26|土地里上好的初熟之物要奉到耶和华－你上帝的殿。不可用母山羊的奶来煮它的小山羊。”
EXOD|34|27|耶和华对 摩西 说：“你要将这些话写上，因为我按这话与你和 以色列 人立约。”
EXOD|34|28|摩西 在耶和华那里四十昼夜，不吃饭不喝水。他把这约的话，那十条诫命 ，写在版上。
EXOD|34|29|摩西 下 西奈山 。 摩西 从山上下来的时候，手里拿着两块法版。 摩西 不知道自己脸上的皮肤因耶和华和他说话而发光。
EXOD|34|30|亚伦 和 以色列 众人看见 摩西 ，看哪，他脸上的皮肤发光，他们就怕靠近他。
EXOD|34|31|摩西 叫他们来， 亚伦 和会众的官长回到他那里， 摩西 就跟他们说话。
EXOD|34|32|随后 以色列 众人都近前来，他就把耶和华在 西奈山 与他所说的一切话都吩咐他们。
EXOD|34|33|摩西 跟他们说完了话，就用面纱蒙上脸。
EXOD|34|34|但 摩西 进到耶和华面前与他说话的时候，就把面纱揭下，直到出来。 摩西 出来，将所吩咐他的话告诉 以色列 人。
EXOD|34|35|以色列 人看见 摩西 的脸，他脸上的皮肤发光。 摩西 就用面纱蒙上脸，直到他进去与耶和华说话才揭下。
EXOD|35|1|摩西 召集 以色列 全会众，对他们说：“这是耶和华吩咐你们遵行的事：
EXOD|35|2|六日要做工，第七日你们要奉为向耶和华守完全安息的安息圣日。凡在这日做工的，要被处死。
EXOD|35|3|在安息日这一天，不可在你们一切的住处生火。”
EXOD|35|4|摩西 对 以色列 全会众说：“这是耶和华所吩咐的话，说：
EXOD|35|5|要从你们当中拿礼物献给耶和华；凡甘心乐意的，可以把耶和华的礼物拿来，就是金、银、铜，
EXOD|35|6|蓝色、紫色、朱红色纱，细麻，山羊毛，
EXOD|35|7|染红的公羊皮，精美的皮料，金合欢木，
EXOD|35|8|点灯的油，做膏油的香料、做香的香料，
EXOD|35|9|红玛瑙与宝石，可以镶嵌在以弗得和胸袋上。”
EXOD|35|10|“你们当中凡心里有智慧的都要来，制造一切耶和华所吩咐的，
EXOD|35|11|就是帐幕、帐幕的罩棚、帐幕的盖、钩子、竖板、横木、柱子和带卯眼的座，
EXOD|35|12|柜子、柜子的杠、柜盖和遮掩的幔子，
EXOD|35|13|供桌、供桌的杠、供桌一切的器具和供饼，
EXOD|35|14|灯台、灯台的器具、灯和点灯的油，
EXOD|35|15|香坛、坛的杠、膏油和芬芳的香，帐幕门口的门帘，
EXOD|35|16|燔祭坛、坛的铜网、坛的杠和坛的一切器具，洗濯盆和盆座，
EXOD|35|17|院子的帷幔、柱子、带卯眼的座和院子的门帘，
EXOD|35|18|帐幕的橛子、院子的橛子和绳子，
EXOD|35|19|以及圣所事奉用的精致礼服， 亚伦 祭司的圣衣和他儿子的衣服，供祭司职分用。”
EXOD|35|20|以色列 全会众从 摩西 的面前出去。
EXOD|35|21|凡心受感动，灵被驱策的，都带耶和华的礼物来，为要造会幕和其中一切的器具，以及缝制圣衣。
EXOD|35|22|凡甘心乐意的，连男带女都来了，各将金器，就是胸针、耳环、打印的戒指，和项链带来，摇着金器的摇祭献给耶和华。
EXOD|35|23|凡有蓝色、紫色、朱红色纱、细麻、山羊毛、染红的公羊皮、精美皮料的，都拿了来；
EXOD|35|24|凡愿意献银和铜作礼物的，都拿礼物来献给耶和华；凡有金合欢木可做各种用途的也都拿了来。
EXOD|35|25|凡心中有智慧，可以亲手纺织的妇女，也把所纺的蓝色、紫色、朱红色纱，和细麻都拿了来。
EXOD|35|26|凡有智慧，心里受感动的妇女都来纺山羊毛。
EXOD|35|27|众官长把红玛瑙和宝石，可以镶嵌在以弗得与胸袋上的，都拿了来，
EXOD|35|28|又拿做香，做膏油，和点灯所需的香料和油来。
EXOD|35|29|以色列 人，无论男女，凡心里受感动的，都带甘心祭来献给耶和华，为要做耶和华藉 摩西 所吩咐的一切工。
EXOD|35|30|摩西 对 以色列 人说：“看， 犹大 支派中 户珥 的孙子， 乌利 的儿子 比撒列 ，耶和华已经题名召他，
EXOD|35|31|又以上帝的灵充满他，使他有智慧、聪明、知识，能做各样的工，
EXOD|35|32|能设计图案，用金、银、铜制造各物，
EXOD|35|33|又能雕刻镶嵌用的宝石，雕刻木头，做各样精巧的工。
EXOD|35|34|耶和华又赐给他和 但 支派中， 亚希撒抹 的儿子 亚何利亚伯 能教导人的心。
EXOD|35|35|耶和华使他们的心满有智慧，能做各样的工，无论是雕刻的工，图案设计的工，用蓝色、紫色、朱红色纱，和细麻作刺绣的工，以及编织的工，他们都能胜任，也能设计图案。”
EXOD|36|1|比撒列 和 亚何利亚伯 ，以及一切心里有智慧，蒙耶和华赐智慧和聪明，懂得做圣所各样用途之工的人，都照耶和华所吩咐的去做。
EXOD|36|2|摩西 把 比撒列 和 亚何利亚伯 ，以及那些蒙耶和华赐他心里有智慧，心受感动愿意前来做工的人都召来。
EXOD|36|3|这些人就从 摩西 收了 以色列 人为建造圣所，以及圣所各用途之工而奉献的礼物。每天早晨，百姓继续把甘心祭拿来。
EXOD|36|4|凡有智慧能做圣所一切工的人，都各自离开他们原本的工作前来，
EXOD|36|5|对 摩西 说：“百姓送来的礼物很多，已经超过耶和华吩咐建造之工所需要的了。”
EXOD|36|6|摩西 吩咐，他们就在营中传令说：“无论男女，不必再为圣所的礼物做任何的工。”这样才使百姓停止，不再拿礼物来，
EXOD|36|7|他们所有的材料已经足够整个工程之用，而且有余。
EXOD|36|8|做工的人当中，凡心里有智慧的，用十幅幔子做帐幕，幔子是用搓的细麻和蓝色、紫色、朱红色纱织成的，并且以刺绣的手艺绣上基路伯。
EXOD|36|9|每幅幔子长二十八肘，每幅幔子宽四肘，全部的幔子都是一样的尺寸。
EXOD|36|10|他使这五幅幔子彼此相连，又使那五幅幔子彼此相连。
EXOD|36|11|他在这一组相连幔子的末幅边上缝了蓝色的钮环；在另一组相连幔子的末幅边上也照样做。
EXOD|36|12|他在这幅幔子上缝五十个钮环，在另一组相连幔子的末幅上也缝五十个钮环，环环相对。
EXOD|36|13|他又做了五十个金钩，用钩子使幔子彼此相连，成为一个帐幕。
EXOD|36|14|他用山羊毛织十一幅幔子，作为帐幕上的罩棚。
EXOD|36|15|每幅幔子长三十肘，每幅幔子宽四肘；十一幅幔子都是一样的尺寸。
EXOD|36|16|他把五幅幔子连成一幅，又把六幅幔子连成一幅。
EXOD|36|17|他在这一组相连幔子的末幅边上缝了五十个钮环；在另一组相连幔子的末幅边上也缝了五十个钮环。
EXOD|36|18|他又做五十个铜钩，使罩棚相连成为一个。
EXOD|36|19|他用染红的公羊皮做罩棚的盖，再用精美皮料做外层的盖。
EXOD|36|20|他用金合欢木做竖立帐幕的木板，
EXOD|36|21|木板长十肘，每块板宽一肘半，
EXOD|36|22|每块板有两个榫头可以彼此衔接。帐幕一切的板都是这样做。
EXOD|36|23|他做帐幕的木板：南面，就是面向南方的那一边，做二十块板，
EXOD|36|24|在这二十块板底下做了四十个带卯眼的银座：两个卯眼接连这块板上的两个榫头，另外两个卯眼接连那块板上的两个榫头。
EXOD|36|25|他在帐幕的第二边，就是北面，也做二十块板，
EXOD|36|26|和四十个带卯眼的银座；这块板底下有两个卯眼，那块板底下也有两个卯眼。
EXOD|36|27|他在帐幕的后面，就是西面，做六块板，
EXOD|36|28|在帐幕后面的角落做两块板。
EXOD|36|29|下端的板是成双的，上端连在一起，直到顶端的第一个环子；两块板都是这样，做成两个角落。
EXOD|36|30|一共有八块板和十六个带卯眼的银座，每块板底下有两个卯眼。
EXOD|36|31|他用金合欢木做横木：为帐幕这面的板做五根横木，
EXOD|36|32|为帐幕那面的板做五根横木，又为帐幕后面，就是朝西的板做五根横木，
EXOD|36|33|他做了板腰间的横木，从一头通到另一头。
EXOD|36|34|他将板包上金子，又做板上的金环来套横木；横木也包上金子。
EXOD|36|35|他用蓝色、紫色、朱红色纱，和搓的细麻织幔子，以刺绣的手艺绣上基路伯。
EXOD|36|36|他又用金合欢木为幔子做四根柱子，包上金子，柱子有金钩，又为柱子铸了四个带卯眼的银座。
EXOD|36|37|他用蓝色、紫色、朱红色纱，和搓的细麻，以刺绣的手艺为帐幕织门帘，
EXOD|36|38|又为帘子做五根柱子和柱子的钩子，把柱顶和柱子的箍包上金子。柱子有五个带卯眼的铜座。
EXOD|37|1|比撒列 用金合欢木做一个柜子，长二肘半，宽一肘半，高一肘半。
EXOD|37|2|里里外外包上金子，四围镶上金边。
EXOD|37|3|他又铸了四个金环，安在柜子的四脚上；这边两个环，那边两个环。
EXOD|37|4|他用金合欢木做了两根杠，包上金子，
EXOD|37|5|又把杠穿过柜旁的环，以便抬柜。
EXOD|37|6|他用纯金做了一个柜盖，长二肘半，宽一肘半，
EXOD|37|7|他造两个用金子锤出的基路伯，从柜盖的两端锤出它们。
EXOD|37|8|这端一个基路伯，那端一个基路伯；从柜盖的两端锤出两个基路伯。
EXOD|37|9|二基路伯的翅膀向上张开，用翅膀遮住柜盖，脸彼此相对；基路伯的脸朝向柜盖。
EXOD|37|10|他用金合欢木做了一张供桌，长二肘，宽一肘，高一肘半，
EXOD|37|11|把它包上纯金，四围镶上金边。
EXOD|37|12|供桌的四围各做了一掌宽的边缘，边缘镶上金边。
EXOD|37|13|他又铸了四个金环，把环安在四个桌脚的四角上。
EXOD|37|14|环靠近边缘，以便穿杠抬供桌。
EXOD|37|15|他用金合欢木做了两根杠，包上金子，用来抬供桌。
EXOD|37|16|他又用纯金做了桌上的器具，就是盘、碟，以及浇酒祭的杯和壶。
EXOD|37|17|他造一座用纯金锤出的灯台；灯台的座、干、杯、花萼和花瓣，都和灯台接连一块。
EXOD|37|18|灯台两旁伸出六根枝子：这边三根，那边三根。
EXOD|37|19|这边的枝子上有三个杯，形状像杏花，有花萼有花瓣；那边的枝子上也有三个杯，形状像杏花，有花萼有花瓣。从灯台伸出来的六根枝子都是如此。
EXOD|37|20|灯台本身有四个杯，形状像杏花，有花萼有花瓣。
EXOD|37|21|灯台的第一对枝子下面有花萼，灯台的第二对枝子下面有花萼，灯台的第三对枝子下面也有花萼；灯台伸出的六根枝子都是如此。
EXOD|37|22|花萼和枝子都和灯台接连一块，全是从一块纯金锤出来的。
EXOD|37|23|他用纯金做灯台的七盏灯，以及灯剪和灯盘。
EXOD|37|24|他用一他连得的纯金做灯台和灯台的一切器具。
EXOD|37|25|他用金合欢木做香坛，长一肘，宽一肘，这坛是正方形的，高二肘。坛的四个翘角与坛接连一块。
EXOD|37|26|他把坛的上面与坛的四围，以及坛的四个翘角包上纯金，又在坛的四围镶上金边。
EXOD|37|27|他在坛的两个对侧，金边下面做了两个金环，用来穿杠抬坛。
EXOD|37|28|他又用金合欢木做杠，包上金子。
EXOD|37|29|他按配制香料的方法制成圣膏油和芬芳的纯香。
EXOD|38|1|他用金合欢木做燔祭坛，长五肘，宽五肘，是正方形的，高三肘。
EXOD|38|2|在坛的四角做四个翘角，与坛接连一块，把坛包上铜。
EXOD|38|3|他做坛的一切器具，就是桶子、铲子、盘子、肉叉和火盆；这一切器具都是用铜做的。
EXOD|38|4|他又为坛做一个铜网，安在坛四围的边的下面，垂到坛的半腰。
EXOD|38|5|他在铜网的四角上铸了四个环，用来穿杠。
EXOD|38|6|他用金合欢木做杠，包上铜，
EXOD|38|7|把杠穿过坛两旁的环子，用来抬坛。他用板做坛，坛的中心是空的。
EXOD|38|8|他用铜做洗濯盆和盆座，是用会幕门前事奉之妇人的铜镜做的。
EXOD|38|9|他又做院子，在南面，就是面向南方的那一边，用搓的细麻做院子的帷幔，一百肘。
EXOD|38|10|帷幔有二十根柱子，二十个带卯眼的铜座；柱子的钩和箍都是银的。
EXOD|38|11|北面的帷幔一百肘。帷幔有二十根柱子，二十个带卯眼的铜座；柱子的钩和箍都是银的。
EXOD|38|12|西面的帷幔五十肘。帷幔有十根柱子，十个带卯眼的座；柱子的钩和箍都是银的。
EXOD|38|13|院子的东面，就是面向东方的那一边，五十肘。
EXOD|38|14|一边的帷幔有十五肘，有三根柱子，三个带卯眼的座。
EXOD|38|15|另一边也一样，院子门口左右的帷幔也有十五肘，有三根柱子，三个带卯眼的座。
EXOD|38|16|院子四面的帷幔都是用搓的细麻做的。
EXOD|38|17|柱子带卯眼的座是铜的，柱子的钩和箍是银的，柱顶是用银包的。院子一切的柱子都是用银子箍着的。
EXOD|38|18|院子的门帘是以刺绣的手艺，用蓝色、紫色、朱红色纱，和搓的细麻织的，长二十肘，宽也就是高五肘，与院子帷幔的高度相同。
EXOD|38|19|门帘有四根柱子，四个带卯眼的铜座；柱子上的钩和箍是银的，柱顶是用银包的。
EXOD|38|20|帐幕一切的橛子和院子四围的橛子都是铜的。
EXOD|38|21|这是帐幕，就是法柜帐幕中物件的总数，是照 摩西 的吩咐， 亚伦 祭司的儿子 以他玛 经手， 利未 人数点的。
EXOD|38|22|凡耶和华吩咐 摩西 的，都是由 犹大 支派中 户珥 的孙子， 乌利 的儿子 比撒列 去做的；
EXOD|38|23|与他同工的有 但 支派中 亚希撒抹 的儿子 亚何利亚伯 ；他是雕刻师，也是设计师，又是用蓝色、紫色、朱红色纱，和细麻的刺绣师。
EXOD|38|24|为圣所一切工作用的金子，就是所奉献的金子，按圣所的舍客勒，一共是二十九他连得，七百三十舍客勒。
EXOD|38|25|会中被数的人所献的银子，按圣所的舍客勒，一共是一百他连得，一千七百七十五舍客勒。
EXOD|38|26|凡曾被数的，就是二十岁以上的人，共有六十万三千五百五十人。按圣所的舍客勒，每人半舍客勒，就是一比加。
EXOD|38|27|一百他连得银子是用来铸造圣所带卯眼的座和幔子下带卯眼的座；用一百他连得铸造一百个带卯眼的座，每个带卯眼的座一他连得。
EXOD|38|28|一千七百七十五舍客勒是用来铸造柱子的钩，包柱顶，以及箍着柱子。
EXOD|38|29|所奉献的铜共有七十他连得，二千四百舍客勒。
EXOD|38|30|这些铜是用来做会幕门口带卯眼的座，铜坛、坛的铜网和坛的一切器具，
EXOD|38|31|院子四围带卯眼的座和院子门口带卯眼的座，以及帐幕一切的橛子和院子四围所有的橛子。
EXOD|39|1|他们用蓝色、紫色、朱红色纱缝制精致的礼服，在圣所用以供职；他们为 亚伦 做圣衣，是照耶和华所吩咐 摩西 的。
EXOD|39|2|以弗得是用金色、蓝色、紫色、朱红色纱，和搓的细麻做的。
EXOD|39|3|他们把金子锤成薄片，剪成细线，与蓝色、紫色、朱红色纱，以刺绣的手艺织在一起。
EXOD|39|4|他们又为以弗得做两条相连的肩带，接连在以弗得的两端。
EXOD|39|5|以弗得的精致带子以一样的手艺，用金色、蓝色、紫色、朱红色纱，和搓的细麻缝制，与以弗得接连在一起，是照耶和华所吩咐 摩西 的。
EXOD|39|6|他们琢出两块红玛瑙，镶在金槽里，如同刻印章，刻上 以色列 众子的名字。
EXOD|39|7|他把这两块宝石安在以弗得的两条肩带上，为 以色列 人作纪念石，是照耶和华所吩咐 摩西 的。
EXOD|39|8|胸袋是以刺绣的手艺，如同以弗得的做法，用金色、蓝色、紫色、朱红色纱，和搓的细麻缝制。
EXOD|39|9|胸袋是正方形的，他们把它做成两层，这两层各长一虎口，宽一虎口。
EXOD|39|10|他们在上面镶四行宝石：第一行是红宝石、红璧玺、红玉；
EXOD|39|11|第二行是绿宝石、蓝宝石、金刚石；
EXOD|39|12|第三行是紫玛瑙、白玛瑙、紫晶；
EXOD|39|13|第四行是水苍玉、红玛瑙、碧玉。这些都镶在金槽中。
EXOD|39|14|这些宝石有 以色列 十二个儿子的名字，如同刻印章，每一颗有自己的名字，代表十二个支派。
EXOD|39|15|他们在胸袋上用纯金打链子，像编成的绳子一样。
EXOD|39|16|他们又做了两个金槽和两个金环，把这两个环安在胸袋的两端。
EXOD|39|17|他们把那两条编成的金链系在胸袋两端的两个环上，
EXOD|39|18|又把链子的另外两端扣在两个槽上，安在以弗得前面的肩带上。
EXOD|39|19|他们做了两个金环，安在胸袋的两端，在以弗得里面的边上，
EXOD|39|20|又做两个金环，安在以弗得前面两条肩带的下边，靠近接缝处，在精致带子的上面。
EXOD|39|21|他们用蓝色的带子把胸袋的环与以弗得的环系住，使胸袋绑在以弗得精致的带子上，不致松脱，是照耶和华所吩咐 摩西 的。
EXOD|39|22|以弗得的外袍是以编织的手艺做的，颜色全是蓝的。
EXOD|39|23|袍上方的中间留了一个领口，领口的周围织出领边，好像铠甲的领口，免得破裂。
EXOD|39|24|他们在袍子下摆用蓝色、紫色、朱红色纱，和搓的细麻 做石榴，
EXOD|39|25|又用纯金铸了铃铛，把铃铛钉在石榴中间，袍子下摆周围的石榴中间：
EXOD|39|26|一个铃铛一个石榴，一个铃铛一个石榴，在袍子下摆的周围，用以供职，是照耶和华所吩咐 摩西 的。
EXOD|39|27|他们用编织的工为 亚伦 和他的儿子做细麻布内袍、
EXOD|39|28|细麻布礼冠、细麻布精致头巾，和搓的细麻布裤子，
EXOD|39|29|又用蓝色、紫色、朱红色纱，和搓的细麻，以刺绣的手艺做腰带，是照耶和华所吩咐 摩西 的。
EXOD|39|30|他们用纯金做一面圣冠上的牌，如同刻印章，在上面写着“归耶和华为圣”，
EXOD|39|31|又用蓝色的带子把牌系在礼冠上，是照耶和华所吩咐 摩西 的。
EXOD|39|32|会幕的帐幕一切的工程就这样做完了。凡耶和华所吩咐 摩西 的， 以色列 人都照样做了。
EXOD|39|33|他们把帐幕运到 摩西 那里，帐幕和帐幕的一切器具，就是钩、板、横木、柱子、带卯眼的座，
EXOD|39|34|染红公羊皮的盖、精美皮料的盖、遮掩的幔子，
EXOD|39|35|法柜、柜的杠、柜盖，
EXOD|39|36|供桌、供桌的一切器具、供饼，
EXOD|39|37|纯金的灯台、摆列的灯、灯台的一切器具、点灯的油，
EXOD|39|38|金坛、膏油、芬芳的香、帐幕的门帘，
EXOD|39|39|铜坛、坛的铜网、坛的杠、坛的一切器具，洗濯盆和盆座，
EXOD|39|40|院子的帷幔、柱子、带卯眼的座、院子的门帘、绳子、橛子，帐幕，就是会幕使用的一切器具，
EXOD|39|41|以及圣所事奉用的精致礼服， 亚伦 祭司的圣衣和他儿子的衣服，供祭司职分用。
EXOD|39|42|这一切工作都是 以色列 人照耶和华所吩咐 摩西 做的。
EXOD|39|43|摩西 看见这一切的工，看哪，耶和华怎样吩咐，他们就照样做了， 摩西 就为他们祝福。
EXOD|40|1|耶和华吩咐 摩西 说：
EXOD|40|2|“正月初一，你要立起会幕的帐幕，
EXOD|40|3|把法柜安放在里面，用幔子将柜遮掩。
EXOD|40|4|把供桌搬进去，摆设桌上的器具。又把灯台搬进去，点上灯。
EXOD|40|5|把金香坛安在法柜前，挂上帐幕的门帘。
EXOD|40|6|把燔祭坛安在会幕的帐幕门前。
EXOD|40|7|把洗濯盆安在会幕和坛的中间，在盆里盛水。
EXOD|40|8|又要在院子周围支起帷幔，把院子的门帘挂上。
EXOD|40|9|你要用膏油抹帐幕和其中所有的，使帐幕和一切器具分别为圣，就都成为圣。
EXOD|40|10|又要抹燔祭坛和坛的一切器具，使坛分别为圣，坛就成为至圣。
EXOD|40|11|要抹洗濯盆和盆座，使盆分别为圣。
EXOD|40|12|你要带 亚伦 和他儿子到会幕门口，用水洗身。
EXOD|40|13|要给 亚伦 穿上圣衣，又膏他，使他分别为圣，作事奉我的祭司。
EXOD|40|14|又要带他的儿子来，给他们穿上内袍。
EXOD|40|15|你怎样膏他们的父亲，也要照样膏他们，使他们成为事奉我的祭司。他们受了膏，就必世世代代永远得祭司的职分。”
EXOD|40|16|摩西 这样做了；耶和华怎样吩咐 摩西 ，他就照样做了。
EXOD|40|17|第二年正月初一，帐幕就立起来。
EXOD|40|18|摩西 支起帐幕，安上带卯眼的座，安上板，穿上横木，立起柱子。
EXOD|40|19|他在帐幕的上面搭上罩棚，把罩棚外层的盖子盖在其上，是照着耶和华所吩咐他的。
EXOD|40|20|他把法版放在柜里，把杠穿在柜的两旁，把柜盖安在柜上。
EXOD|40|21|把柜抬进帐幕，挂上遮掩柜的幔子，把法柜遮盖了，是照耶和华所吩咐 摩西 的。
EXOD|40|22|他把供桌安在会幕内，在帐幕的北边，幔子的外面。
EXOD|40|23|把饼摆设在供桌上，在耶和华面前，是照耶和华所吩咐 摩西 的。
EXOD|40|24|他把灯台安在会幕内，在帐幕的南边，供桌的对面，
EXOD|40|25|并在耶和华面前点灯，是照耶和华所吩咐 摩西 的。
EXOD|40|26|他把金坛安在会幕内，幔子的前面，
EXOD|40|27|又在坛上烧芬芳的香，是照耶和华所吩咐 摩西 的。
EXOD|40|28|他又挂上帐幕的门帘。
EXOD|40|29|在会幕的帐幕门口安设燔祭坛，把燔祭和素祭献在坛上，是照耶和华所吩咐 摩西 的。
EXOD|40|30|他又把洗濯盆安在会幕和祭坛的中间，盆里盛水，以便洗濯。
EXOD|40|31|摩西 和 亚伦 ，以及 亚伦 的儿子用这盆洗手洗脚。
EXOD|40|32|他们进会幕或走近坛的时候，就都洗濯，是照耶和华所吩咐 摩西 的。
EXOD|40|33|他在帐幕和祭坛的四围支起院子的帷幔，把院子的门帘挂上。这样， 摩西 就做完了工。
EXOD|40|34|那时，云彩遮盖会幕，耶和华的荣光充满了帐幕。
EXOD|40|35|摩西 不能进会幕，因为云彩停在其上，耶和华的荣光充满了帐幕。
EXOD|40|36|每逢云彩从帐幕升上去， 以色列 人就起程前行；
EXOD|40|37|云彩若不升上去，他们就不起程，直等到云彩升上去。
EXOD|40|38|在他们所行的路上，在 以色列 全家的眼前，白天，耶和华的云彩在帐幕上，黑夜，有火在云彩中。
