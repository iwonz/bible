ZECH|1|1|In the eighth month of the second year of Darius, the word of the LORD came to the prophet Zechariah son of Berekiah, the son of Iddo:
ZECH|1|2|"The LORD was very angry with your forefathers.
ZECH|1|3|Therefore tell the people: This is what the LORD Almighty says: 'Return to me,' declares the LORD Almighty, 'and I will return to you,' says the LORD Almighty.
ZECH|1|4|Do not be like your forefathers, to whom the earlier prophets proclaimed: This is what the LORD Almighty says: 'Turn from your evil ways and your evil practices.' But they would not listen or pay attention to me, declares the LORD.
ZECH|1|5|Where are your forefathers now? And the prophets, do they live forever?
ZECH|1|6|But did not my words and my decrees, which I commanded my servants the prophets, overtake your forefathers? "Then they repented and said, 'The LORD Almighty has done to us what our ways and practices deserve, just as he determined to do.'" The Man Among the Myrtle Trees
ZECH|1|7|On the twenty-fourth day of the eleventh month, the month of Shebat, in the second year of Darius, the word of the LORD came to the prophet Zechariah son of Berekiah, the son of Iddo.
ZECH|1|8|During the night I had a vision-and there before me was a man riding a red horse! He was standing among the myrtle trees in a ravine. Behind him were red, brown and white horses.
ZECH|1|9|I asked, "What are these, my lord?" The angel who was talking with me answered, "I will show you what they are."
ZECH|1|10|Then the man standing among the myrtle trees explained, "They are the ones the LORD has sent to go throughout the earth."
ZECH|1|11|And they reported to the angel of the LORD, who was standing among the myrtle trees, "We have gone throughout the earth and found the whole world at rest and in peace."
ZECH|1|12|Then the angel of the LORD said, "LORD Almighty, how long will you withhold mercy from Jerusalem and from the towns of Judah, which you have been angry with these seventy years?"
ZECH|1|13|So the LORD spoke kind and comforting words to the angel who talked with me.
ZECH|1|14|Then the angel who was speaking to me said, "Proclaim this word: This is what the LORD Almighty says: 'I am very jealous for Jerusalem and Zion,
ZECH|1|15|but I am very angry with the nations that feel secure. I was only a little angry, but they added to the calamity.'
ZECH|1|16|"Therefore, this is what the LORD says: 'I will return to Jerusalem with mercy, and there my house will be rebuilt. And the measuring line will be stretched out over Jerusalem,' declares the LORD Almighty.
ZECH|1|17|"Proclaim further: This is what the LORD Almighty says: 'My towns will again overflow with prosperity, and the LORD will again comfort Zion and choose Jerusalem.'"
ZECH|1|18|Then I looked up-and there before me were four horns!
ZECH|1|19|I asked the angel who was speaking to me, "What are these?" He answered me, "These are the horns that scattered Judah, Israel and Jerusalem."
ZECH|1|20|Then the LORD showed me four craftsmen.
ZECH|1|21|I asked, "What are these coming to do?" He answered, "These are the horns that scattered Judah so that no one could raise his head, but the craftsmen have come to terrify them and throw down these horns of the nations who lifted up their horns against the land of Judah to scatter its people."
ZECH|2|1|Then I looked up-and there before me was a man with a measuring line in his hand!
ZECH|2|2|I asked, "Where are you going?" He answered me, "To measure Jerusalem, to find out how wide and how long it is."
ZECH|2|3|Then the angel who was speaking to me left, and another angel came to meet him
ZECH|2|4|and said to him: "Run, tell that young man, 'Jerusalem will be a city without walls because of the great number of men and livestock in it.
ZECH|2|5|And I myself will be a wall of fire around it,' declares the LORD, 'and I will be its glory within.'
ZECH|2|6|"Come! Come! Flee from the land of the north," declares the LORD, "for I have scattered you to the four winds of heaven," declares the LORD.
ZECH|2|7|"Come, O Zion! Escape, you who live in the Daughter of Babylon!"
ZECH|2|8|For this is what the LORD Almighty says: "After he has honored me and has sent me against the nations that have plundered you-for whoever touches you touches the apple of his eye-
ZECH|2|9|I will surely raise my hand against them so that their slaves will plunder them. Then you will know that the LORD Almighty has sent me.
ZECH|2|10|"Shout and be glad, O Daughter of Zion. For I am coming, and I will live among you," declares the LORD.
ZECH|2|11|"Many nations will be joined with the LORD in that day and will become my people. I will live among you and you will know that the LORD Almighty has sent me to you.
ZECH|2|12|The LORD will inherit Judah as his portion in the holy land and will again choose Jerusalem.
ZECH|2|13|Be still before the LORD, all mankind, because he has roused himself from his holy dwelling."
ZECH|3|1|Then he showed me Joshua the high priest standing before the angel of the LORD, and Satan standing at his right side to accuse him.
ZECH|3|2|The LORD said to Satan, "The LORD rebuke you, Satan! The LORD, who has chosen Jerusalem, rebuke you! Is not this man a burning stick snatched from the fire?"
ZECH|3|3|Now Joshua was dressed in filthy clothes as he stood before the angel.
ZECH|3|4|The angel said to those who were standing before him, "Take off his filthy clothes." Then he said to Joshua, "See, I have taken away your sin, and I will put rich garments on you."
ZECH|3|5|Then I said, "Put a clean turban on his head." So they put a clean turban on his head and clothed him, while the angel of the LORD stood by.
ZECH|3|6|The angel of the LORD gave this charge to Joshua:
ZECH|3|7|"This is what the LORD Almighty says: 'If you will walk in my ways and keep my requirements, then you will govern my house and have charge of my courts, and I will give you a place among these standing here.
ZECH|3|8|"'Listen, O high priest Joshua and your associates seated before you, who are men symbolic of things to come: I am going to bring my servant, the Branch.
ZECH|3|9|See, the stone I have set in front of Joshua! There are seven eyes on that one stone, and I will engrave an inscription on it,' says the LORD Almighty, 'and I will remove the sin of this land in a single day.
ZECH|3|10|"'In that day each of you will invite his neighbor to sit under his vine and fig tree,' declares the LORD Almighty."
ZECH|4|1|Then the angel who talked with me returned and wakened me, as a man is wakened from his sleep.
ZECH|4|2|He asked me, "What do you see?" I answered, "I see a solid gold lampstand with a bowl at the top and seven lights on it, with seven channels to the lights.
ZECH|4|3|Also there are two olive trees by it, one on the right of the bowl and the other on its left."
ZECH|4|4|I asked the angel who talked with me, "What are these, my lord?"
ZECH|4|5|He answered, "Do you not know what these are?No, my lord," I replied.
ZECH|4|6|So he said to me, "This is the word of the LORD to Zerubbabel: 'Not by might nor by power, but by my Spirit,' says the LORD Almighty.
ZECH|4|7|"What are you, O mighty mountain? Before Zerubbabel you will become level ground. Then he will bring out the capstone to shouts of 'God bless it! God bless it!'"
ZECH|4|8|Then the word of the LORD came to me:
ZECH|4|9|"The hands of Zerubbabel have laid the foundation of this temple; his hands will also complete it. Then you will know that the LORD Almighty has sent me to you.
ZECH|4|10|"Who despises the day of small things? Men will rejoice when they see the plumb line in the hand of Zerubbabel. "(These seven are the eyes of the LORD, which range throughout the earth.)"
ZECH|4|11|Then I asked the angel, "What are these two olive trees on the right and the left of the lampstand?"
ZECH|4|12|Again I asked him, "What are these two olive branches beside the two gold pipes that pour out golden oil?"
ZECH|4|13|He replied, "Do you not know what these are?No, my lord," I said.
ZECH|4|14|So he said, "These are the two who are anointed to serve the Lord of all the earth."
ZECH|5|1|I looked again-and there before me was a flying scroll!
ZECH|5|2|He asked me, "What do you see?" I answered, "I see a flying scroll, thirty feet long and fifteen feet wide. "
ZECH|5|3|And he said to me, "This is the curse that is going out over the whole land; for according to what it says on one side, every thief will be banished, and according to what it says on the other, everyone who swears falsely will be banished.
ZECH|5|4|The LORD Almighty declares, 'I will send it out, and it will enter the house of the thief and the house of him who swears falsely by my name. It will remain in his house and destroy it, both its timbers and its stones.'"
ZECH|5|5|Then the angel who was speaking to me came forward and said to me, "Look up and see what this is that is appearing."
ZECH|5|6|I asked, "What is it?" He replied, "It is a measuring basket. "And he added, "This is the iniquity of the people throughout the land."
ZECH|5|7|Then the cover of lead was raised, and there in the basket sat a woman!
ZECH|5|8|He said, "This is wickedness," and he pushed her back into the basket and pushed the lead cover down over its mouth.
ZECH|5|9|Then I looked up-and there before me were two women, with the wind in their wings! They had wings like those of a stork, and they lifted up the basket between heaven and earth.
ZECH|5|10|"Where are they taking the basket?" I asked the angel who was speaking to me.
ZECH|5|11|He replied, "To the country of Babylonia to build a house for it. When it is ready, the basket will be set there in its place."
ZECH|6|1|I looked up again-and there before me were four chariots coming out from between two mountains-mountains of bronze!
ZECH|6|2|The first chariot had red horses, the second black,
ZECH|6|3|the third white, and the fourth dappled-all of them powerful.
ZECH|6|4|I asked the angel who was speaking to me, "What are these, my lord?"
ZECH|6|5|The angel answered me, "These are the four spirits of heaven, going out from standing in the presence of the Lord of the whole world.
ZECH|6|6|The one with the black horses is going toward the north country, the one with the white horses toward the west, and the one with the dappled horses toward the south."
ZECH|6|7|When the powerful horses went out, they were straining to go throughout the earth. And he said, "Go throughout the earth!" So they went throughout the earth.
ZECH|6|8|Then he called to me, "Look, those going toward the north country have given my Spirit rest in the land of the north."
ZECH|6|9|The word of the LORD came to me:
ZECH|6|10|"Take silver and gold from the exiles Heldai, Tobijah and Jedaiah, who have arrived from Babylon. Go the same day to the house of Josiah son of Zephaniah.
ZECH|6|11|Take the silver and gold and make a crown, and set it on the head of the high priest, Joshua son of Jehozadak.
ZECH|6|12|Tell him this is what the LORD Almighty says: 'Here is the man whose name is the Branch, and he will branch out from his place and build the temple of the LORD.
ZECH|6|13|It is he who will build the temple of the LORD, and he will be clothed with majesty and will sit and rule on his throne. And he will be a priest on his throne. And there will be harmony between the two.'
ZECH|6|14|The crown will be given to Heldai, Tobijah, Jedaiah and Hen son of Zephaniah as a memorial in the temple of the LORD.
ZECH|6|15|Those who are far away will come and help to build the temple of the LORD, and you will know that the LORD Almighty has sent me to you. This will happen if you diligently obey the LORD your God."
ZECH|7|1|In the fourth year of King Darius, the word of the LORD came to Zechariah on the fourth day of the ninth month, the month of Kislev.
ZECH|7|2|The people of Bethel had sent Sharezer and Regem-Melech, together with their men, to entreat the LORD
ZECH|7|3|by asking the priests of the house of the LORD Almighty and the prophets, "Should I mourn and fast in the fifth month, as I have done for so many years?"
ZECH|7|4|Then the word of the LORD Almighty came to me:
ZECH|7|5|"Ask all the people of the land and the priests, 'When you fasted and mourned in the fifth and seventh months for the past seventy years, was it really for me that you fasted?
ZECH|7|6|And when you were eating and drinking, were you not just feasting for yourselves?
ZECH|7|7|Are these not the words the LORD proclaimed through the earlier prophets when Jerusalem and its surrounding towns were at rest and prosperous, and the Negev and the western foothills were settled?'"
ZECH|7|8|And the word of the LORD came again to Zechariah:
ZECH|7|9|"This is what the LORD Almighty says: 'Administer true justice; show mercy and compassion to one another.
ZECH|7|10|Do not oppress the widow or the fatherless, the alien or the poor. In your hearts do not think evil of each other.'
ZECH|7|11|"But they refused to pay attention; stubbornly they turned their backs and stopped up their ears.
ZECH|7|12|They made their hearts as hard as flint and would not listen to the law or to the words that the LORD Almighty had sent by his Spirit through the earlier prophets. So the LORD Almighty was very angry.
ZECH|7|13|"'When I called, they did not listen; so when they called, I would not listen,' says the LORD Almighty.
ZECH|7|14|'I scattered them with a whirlwind among all the nations, where they were strangers. The land was left so desolate behind them that no one could come or go. This is how they made the pleasant land desolate.'"
ZECH|8|1|Again the word of the LORD Almighty came to me.
ZECH|8|2|This is what the LORD Almighty says: "I am very jealous for Zion; I am burning with jealousy for her."
ZECH|8|3|This is what the LORD says: "I will return to Zion and dwell in Jerusalem. Then Jerusalem will be called the City of Truth, and the mountain of the LORD Almighty will be called the Holy Mountain."
ZECH|8|4|This is what the LORD Almighty says: "Once again men and women of ripe old age will sit in the streets of Jerusalem, each with cane in hand because of his age.
ZECH|8|5|The city streets will be filled with boys and girls playing there."
ZECH|8|6|This is what the LORD Almighty says: "It may seem marvelous to the remnant of this people at that time, but will it seem marvelous to me?" declares the LORD Almighty.
ZECH|8|7|This is what the LORD Almighty says: "I will save my people from the countries of the east and the west.
ZECH|8|8|I will bring them back to live in Jerusalem; they will be my people, and I will be faithful and righteous to them as their God."
ZECH|8|9|This is what the LORD Almighty says: "You who now hear these words spoken by the prophets who were there when the foundation was laid for the house of the LORD Almighty, let your hands be strong so that the temple may be built.
ZECH|8|10|Before that time there were no wages for man or beast. No one could go about his business safely because of his enemy, for I had turned every man against his neighbor.
ZECH|8|11|But now I will not deal with the remnant of this people as I did in the past," declares the LORD Almighty.
ZECH|8|12|"The seed will grow well, the vine will yield its fruit, the ground will produce its crops, and the heavens will drop their dew. I will give all these things as an inheritance to the remnant of this people.
ZECH|8|13|As you have been an object of cursing among the nations, O Judah and Israel, so will I save you, and you will be a blessing. Do not be afraid, but let your hands be strong."
ZECH|8|14|This is what the LORD Almighty says: "Just as I had determined to bring disaster upon you and showed no pity when your fathers angered me," says the LORD Almighty,
ZECH|8|15|"so now I have determined to do good again to Jerusalem and Judah. Do not be afraid.
ZECH|8|16|These are the things you are to do: Speak the truth to each other, and render true and sound judgment in your courts;
ZECH|8|17|do not plot evil against your neighbor, and do not love to swear falsely. I hate all this," declares the LORD.
ZECH|8|18|Again the word of the LORD Almighty came to me.
ZECH|8|19|This is what the LORD Almighty says: "The fasts of the fourth, fifth, seventh and tenth months will become joyful and glad occasions and happy festivals for Judah. Therefore love truth and peace."
ZECH|8|20|This is what the LORD Almighty says: "Many peoples and the inhabitants of many cities will yet come,
ZECH|8|21|and the inhabitants of one city will go to another and say, 'Let us go at once to entreat the LORD and seek the LORD Almighty. I myself am going.'
ZECH|8|22|And many peoples and powerful nations will come to Jerusalem to seek the LORD Almighty and to entreat him."
ZECH|8|23|This is what the LORD Almighty says: "In those days ten men from all languages and nations will take firm hold of one Jew by the hem of his robe and say, 'Let us go with you, because we have heard that God is with you.'"
ZECH|9|1|The word of the LORD is against the land of Hadrach and will rest upon Damascus- for the eyes of men and all the tribes of Israel are on the LORD -
ZECH|9|2|and upon Hamath too, which borders on it, and upon Tyre and Sidon, though they are very skillful.
ZECH|9|3|Tyre has built herself a stronghold; she has heaped up silver like dust, and gold like the dirt of the streets.
ZECH|9|4|But the Lord will take away her possessions and destroy her power on the sea, and she will be consumed by fire.
ZECH|9|5|Ashkelon will see it and fear; Gaza will writhe in agony, and Ekron too, for her hope will wither. Gaza will lose her king and Ashkelon will be deserted.
ZECH|9|6|Foreigners will occupy Ashdod, and I will cut off the pride of the Philistines.
ZECH|9|7|I will take the blood from their mouths, the forbidden food from between their teeth. Those who are left will belong to our God and become leaders in Judah, and Ekron will be like the Jebusites.
ZECH|9|8|But I will defend my house against marauding forces. Never again will an oppressor overrun my people, for now I am keeping watch.
ZECH|9|9|Rejoice greatly, O Daughter of Zion! Shout, Daughter of Jerusalem! See, your king comes to you, righteous and having salvation, gentle and riding on a donkey, on a colt, the foal of a donkey.
ZECH|9|10|I will take away the chariots from Ephraim and the war-horses from Jerusalem, and the battle bow will be broken. He will proclaim peace to the nations. His rule will extend from sea to sea and from the River to the ends of the earth.
ZECH|9|11|As for you, because of the blood of my covenant with you, I will free your prisoners from the waterless pit.
ZECH|9|12|Return to your fortress, O prisoners of hope; even now I announce that I will restore twice as much to you.
ZECH|9|13|I will bend Judah as I bend my bow and fill it with Ephraim. I will rouse your sons, O Zion, against your sons, O Greece, and make you like a warrior's sword.
ZECH|9|14|Then the LORD will appear over them; his arrow will flash like lightning. The Sovereign LORD will sound the trumpet; he will march in the storms of the south,
ZECH|9|15|and the LORD Almighty will shield them. They will destroy and overcome with slingstones. They will drink and roar as with wine; they will be full like a bowl used for sprinkling the corners of the altar.
ZECH|9|16|The LORD their God will save them on that day as the flock of his people. They will sparkle in his land like jewels in a crown.
ZECH|9|17|How attractive and beautiful they will be! Grain will make the young men thrive, and new wine the young women.
ZECH|10|1|Ask the LORD for rain in the springtime; it is the LORD who makes the storm clouds. He gives showers of rain to men, and plants of the field to everyone.
ZECH|10|2|The idols speak deceit, diviners see visions that lie; they tell dreams that are false, they give comfort in vain. Therefore the people wander like sheep oppressed for lack of a shepherd.
ZECH|10|3|"My anger burns against the shepherds, and I will punish the leaders; for the LORD Almighty will care for his flock, the house of Judah, and make them like a proud horse in battle.
ZECH|10|4|From Judah will come the cornerstone, from him the tent peg, from him the battle bow, from him every ruler.
ZECH|10|5|Together they will be like mighty men trampling the muddy streets in battle. Because the LORD is with them, they will fight and overthrow the horsemen.
ZECH|10|6|"I will strengthen the house of Judah and save the house of Joseph. I will restore them because I have compassion on them. They will be as though I had not rejected them, for I am the LORD their God and I will answer them.
ZECH|10|7|The Ephraimites will become like mighty men, and their hearts will be glad as with wine. Their children will see it and be joyful; their hearts will rejoice in the LORD.
ZECH|10|8|I will signal for them and gather them in. Surely I will redeem them; they will be as numerous as before.
ZECH|10|9|Though I scatter them among the peoples, yet in distant lands they will remember me. They and their children will survive, and they will return.
ZECH|10|10|I will bring them back from Egypt and gather them from Assyria. I will bring them to Gilead and Lebanon, and there will not be room enough for them.
ZECH|10|11|They will pass through the sea of trouble; the surging sea will be subdued and all the depths of the Nile will dry up. Assyria's pride will be brought down and Egypt's scepter will pass away.
ZECH|10|12|I will strengthen them in the LORD and in his name they will walk," declares the LORD.
ZECH|11|1|Open your doors, O Lebanon, so that fire may devour your cedars!
ZECH|11|2|Wail, O pine tree, for the cedar has fallen; the stately trees are ruined! Wail, oaks of Bashan; the dense forest has been cut down!
ZECH|11|3|Listen to the wail of the shepherds; their rich pastures are destroyed! Listen to the roar of the lions; the lush thicket of the Jordan is ruined!
ZECH|11|4|This is what the LORD my God says: "Pasture the flock marked for slaughter.
ZECH|11|5|Their buyers slaughter them and go unpunished. Those who sell them say, 'Praise the LORD, I am rich!' Their own shepherds do not spare them.
ZECH|11|6|For I will no longer have pity on the people of the land," declares the LORD. "I will hand everyone over to his neighbor and his king. They will oppress the land, and I will not rescue them from their hands."
ZECH|11|7|So I pastured the flock marked for slaughter, particularly the oppressed of the flock. Then I took two staffs and called one Favor and the other Union, and I pastured the flock.
ZECH|11|8|In one month I got rid of the three shepherds. The flock detested me, and I grew weary of them
ZECH|11|9|and said, "I will not be your shepherd. Let the dying die, and the perishing perish. Let those who are left eat one another's flesh."
ZECH|11|10|Then I took my staff called Favor and broke it, revoking the covenant I had made with all the nations.
ZECH|11|11|It was revoked on that day, and so the afflicted of the flock who were watching me knew it was the word of the LORD.
ZECH|11|12|I told them, "If you think it best, give me my pay; but if not, keep it." So they paid me thirty pieces of silver.
ZECH|11|13|And the LORD said to me, "Throw it to the potter"-the handsome price at which they priced me! So I took the thirty pieces of silver and threw them into the house of the LORD to the potter.
ZECH|11|14|Then I broke my second staff called Union, breaking the brotherhood between Judah and Israel.
ZECH|11|15|Then the LORD said to me, "Take again the equipment of a foolish shepherd.
ZECH|11|16|For I am going to raise up a shepherd over the land who will not care for the lost, or seek the young, or heal the injured, or feed the healthy, but will eat the meat of the choice sheep, tearing off their hoofs.
ZECH|11|17|"Woe to the worthless shepherd, who deserts the flock! May the sword strike his arm and his right eye! May his arm be completely withered, his right eye totally blinded!"
ZECH|12|1|This is the word of the LORD concerning Israel. The LORD, who stretches out the heavens, who lays the foundation of the earth, and who forms the spirit of man within him, declares:
ZECH|12|2|"I am going to make Jerusalem a cup that sends all the surrounding peoples reeling. Judah will be besieged as well as Jerusalem.
ZECH|12|3|On that day, when all the nations of the earth are gathered against her, I will make Jerusalem an immovable rock for all the nations. All who try to move it will injure themselves.
ZECH|12|4|On that day I will strike every horse with panic and its rider with madness," declares the LORD. "I will keep a watchful eye over the house of Judah, but I will blind all the horses of the nations.
ZECH|12|5|Then the leaders of Judah will say in their hearts, 'The people of Jerusalem are strong, because the LORD Almighty is their God.'
ZECH|12|6|"On that day I will make the leaders of Judah like a firepot in a woodpile, like a flaming torch among sheaves. They will consume right and left all the surrounding peoples, but Jerusalem will remain intact in her place.
ZECH|12|7|"The LORD will save the dwellings of Judah first, so that the honor of the house of David and of Jerusalem's inhabitants may not be greater than that of Judah.
ZECH|12|8|On that day the LORD will shield those who live in Jerusalem, so that the feeblest among them will be like David, and the house of David will be like God, like the Angel of the LORD going before them.
ZECH|12|9|On that day I will set out to destroy all the nations that attack Jerusalem.
ZECH|12|10|"And I will pour out on the house of David and the inhabitants of Jerusalem a spirit of grace and supplication. They will look on me, the one they have pierced, and they will mourn for him as one mourns for an only child, and grieve bitterly for him as one grieves for a firstborn son.
ZECH|12|11|On that day the weeping in Jerusalem will be great, like the weeping of Hadad Rimmon in the plain of Megiddo.
ZECH|12|12|The land will mourn, each clan by itself, with their wives by themselves: the clan of the house of David and their wives, the clan of the house of Nathan and their wives,
ZECH|12|13|the clan of the house of Levi and their wives, the clan of Shimei and their wives,
ZECH|12|14|and all the rest of the clans and their wives.
ZECH|13|1|"On that day a fountain will be opened to the house of David and the inhabitants of Jerusalem, to cleanse them from sin and impurity.
ZECH|13|2|"On that day, I will banish the names of the idols from the land, and they will be remembered no more," declares the LORD Almighty. "I will remove both the prophets and the spirit of impurity from the land.
ZECH|13|3|And if anyone still prophesies, his father and mother, to whom he was born, will say to him, 'You must die, because you have told lies in the LORD's name.' When he prophesies, his own parents will stab him.
ZECH|13|4|"On that day every prophet will be ashamed of his prophetic vision. He will not put on a prophet's garment of hair in order to deceive.
ZECH|13|5|He will say, 'I am not a prophet. I am a farmer; the land has been my livelihood since my youth. '
ZECH|13|6|If someone asks him, 'What are these wounds on your body?' he will answer, 'The wounds I was given at the house of my friends.'
ZECH|13|7|"Awake, O sword, against my shepherd, against the man who is close to me!" declares the LORD Almighty. "Strike the shepherd, and the sheep will be scattered, and I will turn my hand against the little ones.
ZECH|13|8|In the whole land," declares the LORD, "two-thirds will be struck down and perish; yet one-third will be left in it.
ZECH|13|9|This third I will bring into the fire; I will refine them like silver and test them like gold. They will call on my name and I will answer them; I will say, 'They are my people,' and they will say, 'The LORD is our God.'"
ZECH|14|1|A day of the LORD is coming when your plunder will be divided among you.
ZECH|14|2|I will gather all the nations to Jerusalem to fight against it; the city will be captured, the houses ransacked, and the women raped. Half of the city will go into exile, but the rest of the people will not be taken from the city.
ZECH|14|3|Then the LORD will go out and fight against those nations, as he fights in the day of battle.
ZECH|14|4|On that day his feet will stand on the Mount of Olives, east of Jerusalem, and the Mount of Olives will be split in two from east to west, forming a great valley, with half of the mountain moving north and half moving south.
ZECH|14|5|You will flee by my mountain valley, for it will extend to Azel. You will flee as you fled from the earthquake in the days of Uzziah king of Judah. Then the LORD my God will come, and all the holy ones with him.
ZECH|14|6|On that day there will be no light, no cold or frost.
ZECH|14|7|It will be a unique day, without daytime or nighttime-a day known to the LORD. When evening comes, there will be light.
ZECH|14|8|On that day living water will flow out from Jerusalem, half to the eastern sea and half to the western sea, in summer and in winter.
ZECH|14|9|The LORD will be king over the whole earth. On that day there will be one LORD, and his name the only name.
ZECH|14|10|The whole land, from Geba to Rimmon, south of Jerusalem, will become like the Arabah. But Jerusalem will be raised up and remain in its place, from the Benjamin Gate to the site of the First Gate, to the Corner Gate, and from the Tower of Hananel to the royal winepresses.
ZECH|14|11|It will be inhabited; never again will it be destroyed. Jerusalem will be secure.
ZECH|14|12|This is the plague with which the LORD will strike all the nations that fought against Jerusalem: Their flesh will rot while they are still standing on their feet, their eyes will rot in their sockets, and their tongues will rot in their mouths.
ZECH|14|13|On that day men will be stricken by the LORD with great panic. Each man will seize the hand of another, and they will attack each other.
ZECH|14|14|Judah too will fight at Jerusalem. The wealth of all the surrounding nations will be collected-great quantities of gold and silver and clothing.
ZECH|14|15|A similar plague will strike the horses and mules, the camels and donkeys, and all the animals in those camps.
ZECH|14|16|Then the survivors from all the nations that have attacked Jerusalem will go up year after year to worship the King, the LORD Almighty, and to celebrate the Feast of Tabernacles.
ZECH|14|17|If any of the peoples of the earth do not go up to Jerusalem to worship the King, the LORD Almighty, they will have no rain.
ZECH|14|18|If the Egyptian people do not go up and take part, they will have no rain. The LORD will bring on them the plague he inflicts on the nations that do not go up to celebrate the Feast of Tabernacles.
ZECH|14|19|This will be the punishment of Egypt and the punishment of all the nations that do not go up to celebrate the Feast of Tabernacles.
ZECH|14|20|On that dayHOLY TO THE LORD will be inscribed on the bells of the horses, and the cooking pots in the LORD's house will be like the sacred bowls in front of the altar.
ZECH|14|21|Every pot in Jerusalem and Judah will be holy to the LORD Almighty, and all who come to sacrifice will take some of the pots and cook in them. And on that day there will no longer be a Canaanite in the house of the LORD Almighty.
