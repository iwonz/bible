AMOS|1|1|这是 犹大 王 乌西雅 在位与 约阿施 的儿子 以色列 王 耶罗波安 在位的时候，大地震前二年，从 提哥亚 来的牧人 阿摩司 所见的─他的话论到 以色列 。
AMOS|1|2|他说：“耶和华必从 锡安 吼叫， 从 耶路撒冷 出声； 牧人的草场哀伤， 迦密 的山顶枯干。”
AMOS|1|3|耶和华如此说： “ 大马士革 三番四次犯罪， 以铁的打谷机击打 基列 ， 我必不撤销对它的惩罚。
AMOS|1|4|我要降火在 哈薛 的王宫， 吞灭 便．哈达 的宫殿；
AMOS|1|5|我要折断 大马士革 的门闩， 剪除 亚文 平原的居民 和 伯．伊甸 的掌权者， 亚兰 人必被掳到 吉珥 。” 这是耶和华说的。
AMOS|1|6|耶和华如此说： “ 迦萨 三番四次犯罪， 掳掠全体百姓交给 以东 ， 我必不撤销对它的惩罚。
AMOS|1|7|我要降火在 迦萨 城内， 吞灭它的宫殿；
AMOS|1|8|我要剪除 亚实突 的居民 和 亚实基伦 的掌权者， 反手攻击 以革伦 ， 剩余的 非利士 人都必灭亡。” 这是主耶和华说的。
AMOS|1|9|耶和华如此说： “ 推罗 三番四次犯罪， 将全体百姓交给 以东 ， 不顾念弟兄的盟约， 我必不撤销对它的惩罚，
AMOS|1|10|我要降火在 推罗 城内， 吞灭它的宫殿。”
AMOS|1|11|耶和华如此说： “ 以东 三番四次犯罪， 怒气不停发作，永远怀着愤怒， 拿刀追赶兄弟，丝毫不存怜悯， 我必不撤销对它的惩罚。
AMOS|1|12|我要降火在 提幔 ， 吞灭 波斯拉 的宫殿。”
AMOS|1|13|耶和华如此说： “ 亚扪 人三番四次犯罪， 剖开 基列 的孕妇， 扩张自己的疆界， 我必不撤销对它的惩罚。
AMOS|1|14|我要在战争呐喊的日子， 在旋风狂吹时， 在 拉巴 城内放火， 吞灭它的宫殿；
AMOS|1|15|他们的君王和官长必一同被掳。” 这是耶和华说的。
AMOS|2|1|耶和华如此说： “ 摩押 三番四次犯罪， 把 以东 王的骸骨焚烧成灰， 我必不撤销对它的惩罚。
AMOS|2|2|我要降火在 摩押 ， 吞灭 加略 的宫殿， 摩押 必在闹哄、呐喊、吹角声中灭亡；
AMOS|2|3|我要剪除 摩押 的领袖， 把所有的官长和他一同杀戮。” 这是耶和华说的。
AMOS|2|4|耶和华如此说： “ 犹大 三番四次犯罪， 厌弃耶和华的训诲， 不遵守他的律例； 他们祖先所随从虚假的偶像 使他们走迷了， 我必不撤销对它的惩罚。
AMOS|2|5|我要降火在 犹大 ， 吞灭 耶路撒冷 的宫殿。”
AMOS|2|6|耶和华如此说： “ 以色列 三番四次犯罪， 为银子卖了义人， 为一双鞋卖了穷人， 我必不撤销对它的惩罚。
AMOS|2|7|他们把贫寒人的头践踏在地的尘土上 ， 又阻碍困苦人的道路。 父子与同一个女子行淫， 以致亵渎我的圣名。
AMOS|2|8|他们在各祭坛旁边， 躺卧在人所典当的衣服上， 又在他们上帝的殿里 喝受罚之人的酒。
AMOS|2|9|“我从他们面前除灭 亚摩利 人； 他虽高大如香柏树，强壮如橡树， 我却上灭其果，下绝其根。
AMOS|2|10|我曾将你们从 埃及 地领上来， 在旷野里引导你们四十年， 使你们得 亚摩利 人之地为业；
AMOS|2|11|我从你们子孙中兴起先知， 又从你们少年中兴起拿细耳人。 以色列 人哪，不是这样吗？” 这是耶和华说的。
AMOS|2|12|“你们却把酒给拿细耳人喝， 嘱咐先知说：‘不要说预言。’
AMOS|2|13|“看哪，我要把你们压下去， 如同装满禾捆的车压过一样。
AMOS|2|14|快跑的无从避难， 壮士无法使力， 勇士也不能自救；
AMOS|2|15|拿弓的站立不住， 腿快的不能逃脱， 骑马的也不能自救。
AMOS|2|16|到那日，勇士中最有胆量的， 必赤身逃跑。” 这是耶和华说的。
AMOS|3|1|以色列 人哪，当听耶和华责备你们的话，责备我从 埃及 地领上来的全家，说：
AMOS|3|2|“在地上万族中，我只认识你们； 因此，我必惩罚你们一切的罪孽。”
AMOS|3|3|二人若不同心， 岂能同行呢？
AMOS|3|4|狮子若无猎物， 岂会在林中咆哮呢？ 少壮狮子若无所得， 岂会从洞里吼叫呢？
AMOS|3|5|若未设圈套， 雀鸟岂能陷入地上的罗网呢？ 罗网若无所得， 岂会从地上翻起呢？
AMOS|3|6|城中若吹角， 百姓岂不战兢吗？ 灾祸若临到一城， 岂非耶和华所降的吗？
AMOS|3|7|主耶和华不会做任何事情， 除非先将奥秘指示他的仆人众先知。
AMOS|3|8|狮子吼叫，谁不惧怕呢？ 主耶和华既已说了，谁能不说预言呢？
AMOS|3|9|你们要在 亚实突 的宫殿 和 埃及 地的宫殿传扬，说： “要聚集在 撒玛利亚 的山上， 看城里有何等大的扰乱与欺压。”
AMOS|3|10|“他们以暴力抢夺， 堆积在自己的宫殿里， 却不懂得行正直的事。” 这是耶和华说的。
AMOS|3|11|所以主耶和华如此说： “敌人必来围攻这地， 削弱你的势力， 抢掠你的宫殿。”
AMOS|3|12|耶和华如此说：“牧人怎样从狮子口中抢回两条腿或耳朵的一小片，住 撒玛利亚 的 以色列 人得救也是如此，不过抢回床的一角和床榻的靠枕 而已。”
AMOS|3|13|主耶和华－万军之上帝说： “当听这话，警戒 雅各 家。
AMOS|3|14|我惩罚 以色列 罪孽的日子， 也要惩罚 伯特利 的祭坛； 祭坛的角必被砍下，坠落于地。
AMOS|3|15|我要拆毁过冬和避暑的房屋， 象牙的房屋必毁灭， 广厦豪宅都归无有。” 这是耶和华说的。
AMOS|4|1|“你们这些 撒玛利亚山 上的 巴珊 母牛啊， 当听这话！ 你们欺负贫寒人，压碎贫穷人， 对主人说：‘拿酒来，我们喝吧！’
AMOS|4|2|主耶和华指着自己的神圣起誓说： ‘看哪，日子将到，人必用钩子将你们钩去， 用鱼钩把你们中最后一个钩去。
AMOS|4|3|你们必从城墙的缺口 出去， 各人直往前行， 投向 哈门 。’” 这是耶和华说的。
AMOS|4|4|“ 以色列 人哪，任你们往 伯特利 去犯罪， 到 吉甲 增加罪过， 每早晨献上你们的祭物， 每三日纳你们的十一奉献；
AMOS|4|5|任你们献上有酵的感谢祭， 宣扬你们的甘心祭，使人听见， 因为这是你们所喜爱的。” 这是主耶和华说的。
AMOS|4|6|“我使你们在每一座城里牙齿干净， 使你们各处的粮食缺乏， 你们仍不归向我。” 这是耶和华说的。
AMOS|4|7|“在收割的前三个月， 我不降雨在你们那里， 我降雨在这城， 不降雨在那城； 这块地有雨， 那块无雨的地就必枯干。
AMOS|4|8|两三城的人挤到一个城去找水喝， 却喝不足， 你们仍不归向我。” 这是耶和华说的。
AMOS|4|9|“我以焚风 和霉烂攻击你们， 你们许多的菜园、葡萄园、 无花果树、橄榄树屡屡被剪虫 所吃， 你们仍不归向我。” 这是耶和华说的。
AMOS|4|10|“我降瘟疫在你们中间， 如在 埃及 的样子； 用刀杀戮你们的年轻人 和你们遭掳掠的马匹， 营中臭气扑鼻， 你们仍不归向我。” 这是耶和华说的。
AMOS|4|11|“我倾覆你们， 如同上帝从前倾覆 所多玛 、 蛾摩拉 一样； 你们好像从火中抢救出来的一根柴， 你们仍不归向我。” 这是耶和华说的。
AMOS|4|12|“因此， 以色列 啊，我要如此对待你； 因为我要这样对待你， 以色列 啊， 你当预备迎见你的上帝。”
AMOS|4|13|看哪，那创山，造风，将其心意指示人， 使晨光变幽暗，踩行在地之高处的， 他的名是耶和华－万军之上帝。
AMOS|5|1|以色列 家啊，听我为你们所作的哀歌：
AMOS|5|2|“ 以色列 民 跌倒，不得再起； 躺在地上，无人扶起。”
AMOS|5|3|主耶和华如此说： “ 以色列 家的城派出一千，只剩一百； 派出一百，只剩十个。”
AMOS|5|4|耶和华向 以色列 家如此说： “你们要寻求我，就必存活。
AMOS|5|5|不要往 伯特利 寻求， 不要进入 吉甲 ， 也不要过到 别是巴 ； 因为 吉甲 必被掳走， 伯特利 必归无有。”
AMOS|5|6|要寻求耶和华，就必存活， 免得他在 约瑟 家如火发出， 焚烧 伯特利 ，无人扑灭。
AMOS|5|7|你们这使公平变为茵蔯， 将公义丢弃于地的人哪！
AMOS|5|8|那造昴星和参星， 使死荫变为晨光， 使白昼变为黑夜， 召唤海水、 使其倾倒在地面上的， 耶和华是他的名。
AMOS|5|9|他快速摧毁强壮的人， 毁灭就临到堡垒。
AMOS|5|10|你们怨恨那在城门口断是非的， 憎恶那说正直话的。
AMOS|5|11|所以，因你们践踏贫寒人， 向他们勒索粮税； 你们虽建造石凿的房屋， 却不得住在其内； 虽栽植美好的葡萄园， 却不得喝其中所出的酒。
AMOS|5|12|我知道你们的罪过何其多， 你们的罪恶何其大； 你们迫害义人，收受贿赂， 在城门口屈枉贫穷人。
AMOS|5|13|所以智慧人在这样的时候必静默不言， 因为这是险恶的时候。
AMOS|5|14|你们要寻求良善， 不要寻求邪恶，就必存活。 这样，耶和华－万军之上帝 必照你们所说的与你们同在。
AMOS|5|15|要恨恶邪恶，喜爱良善， 在城门口秉公行义； 或者耶和华－万军之上帝 会施恩给 约瑟 的余民。
AMOS|5|16|因此，主耶和华－万军之上帝如此说： “在一切的广场上必有哀号的声音； 在各街市上必有人说： ‘哀哉！哀哉！’ 他们叫农夫来哭号， 叫善唱哀歌的来举哀；
AMOS|5|17|各葡萄园都有哀号的声音， 因为我必从你中间经过。” 这是耶和华说的。
AMOS|5|18|想望耶和华日子的人有祸了！ 为什么你们要耶和华的日子呢？ 那是黑暗没有光明的日子，
AMOS|5|19|好像人躲避狮子却遇见熊； 进房屋以手靠墙，却被蛇咬。
AMOS|5|20|耶和华的日子岂不是黑暗没有光明， 幽暗毫无光辉吗？
AMOS|5|21|“我厌恶你们的节期， 也不喜悦你们的严肃会。
AMOS|5|22|你们虽然向我献燔祭和素祭， 我却不悦纳， 也不看你们用肥畜献的平安祭。
AMOS|5|23|要使你们歌唱的声音远离我， 因为我不听你们琴瑟的乐曲。
AMOS|5|24|惟愿公平如大水滚滚， 公义如江河滔滔。
AMOS|5|25|“ 以色列 家啊，你们在旷野四十年，何尝将祭物和供物献给我呢？
AMOS|5|26|你们抬着你们的 撒古特 君王 ，和你们为自己所造之偶像 迦温 ，你们的神明之星。
AMOS|5|27|所以我要把你们掳到 大马士革 以外。”这是耶和华说的，他的名为万军之上帝。
AMOS|6|1|“那在 锡安 安逸， 在 撒玛利亚山 安稳， 为列国之首，具有名望， 且为 以色列 家所归向的，有祸了！
AMOS|6|2|你们要过到 甲尼 察看， 从那里往 哈马 大城去， 又下到 非利士 人的 迦特 ， 你们比这些国更好吗？ 或是他们的疆界比你们的疆界广大呢？
AMOS|6|3|你们以为降祸的日子尚远， 却使残暴的统治 临近。
AMOS|6|4|“那些躺卧在象牙床上，舒身在榻上的， 吃群中的羔羊和棚里的牛犊。
AMOS|6|5|他们以琴瑟逍遥歌唱， 为自己作曲 ，像 大卫 一样；
AMOS|6|6|以大碗喝酒，用上等油抹身， 却不为 约瑟 所受的苦难忧伤；
AMOS|6|7|所以，现在这些人必首先被掳， 逍遥的欢宴必消失。”
AMOS|6|8|主耶和华指着自己起誓说： “我憎恶 雅各 的骄傲，厌弃他的宫殿； 我必将城和其中一切所有的都交给敌人。” 这是耶和华－万军之上帝说的 。
AMOS|6|9|那时，若一房之内剩下十个人，也都必死。
AMOS|6|10|死人的叔伯要把尸首抬到屋外焚烧，就问房屋内间的人说：“你那里还有别人吗？”他说：“没有。”又说：“不要作声，不可提耶和华的名。”
AMOS|6|11|看哪，耶和华发命令， 把大房子拆成碎片， 小屋子裂为小块。
AMOS|6|12|马岂能在岩石上奔跑？ 人岂能在那里 用牛耕种呢？ 你们却使公平变为苦胆， 使公义的果子变为茵蔯。
AMOS|6|13|你们这些喜爱 罗．底巴 的，自夸说： “我们不是凭自己的力量攻占了 加宁 吗？”
AMOS|6|14|耶和华─万军之上帝说： “ 以色列 家，看哪，我必兴起一国攻击你们； 他们必欺压你们， 从 哈马口 直到 亚拉巴 的河。”
AMOS|7|1|主耶和华指示我一件事，在春天作物刚长出时，看哪，主 造了蝗虫；看哪，这是王收割后长出的春天作物。
AMOS|7|2|蝗虫吃尽那地青草的时候，我说： “主耶和华啊，求你赦免； 因为 雅各 弱小， 他怎能站立得住呢？”
AMOS|7|3|耶和华对这事改变心意， 耶和华说：“这灾可以免了。”
AMOS|7|4|主耶和华又指示我一件事，看哪，主耶和华命火施行审判，火就吞灭深渊，烧尽产业。
AMOS|7|5|我就说： “主耶和华啊，求你止息； 因为 雅各 弱小， 他怎能站立得住呢？”
AMOS|7|6|耶和华对这事改变心意， 主耶和华说：“这灾也可免了。”
AMOS|7|7|他又指示我一件事，看哪，主手拿铅垂线，站立在依铅垂线建好的墙边。
AMOS|7|8|耶和华对我说：“ 阿摩司 ，你看见什么？”我说：“铅垂线。”主说： “看哪，我要在我子民 以色列 中 吊起铅垂线， 不再宽恕他们。
AMOS|7|9|以撒 的丘坛必荒凉， 以色列 的圣所必荒废； 我要起来用刀攻击 耶罗波安 的家。”
AMOS|7|10|伯特利 的祭司 亚玛谢 派人到 以色列 王 耶罗波安 那里，说：“ 阿摩司 在 以色列 家中图谋背叛你，他所说的一切话，这地不能承担；
AMOS|7|11|因为 阿摩司 这样说： ‘ 耶罗波安 必被刀杀， 以色列 百姓必被掳， 离开本地。’”
AMOS|7|12|于是 亚玛谢 对 阿摩司 说：“你这先见哪，要逃到 犹大 地，在那里过活 ，在那里说预言；
AMOS|7|13|却不要在 伯特利 再说预言，因为这里有王的圣所，有王的宫殿。”
AMOS|7|14|阿摩司 对 亚玛谢 说：“我原不是先知，也不是先知的门徒；我是牧人，是修剪桑树的。
AMOS|7|15|耶和华带领我，叫我不再牧放羊群，对我说：‘你去向我子民 以色列 说预言。’
AMOS|7|16|“现在你要听耶和华的话。 你说：‘不要向 以色列 说预言， 也不要向 以撒 家传讲 。’
AMOS|7|17|所以耶和华如此说： ‘你的妻子要在城中作妓女， 你的儿女要倒在刀下； 你的地必有人用绳子量了瓜分， 你自己必死在不洁净之地； 以色列 百姓必被掳， 离开本地。’”
AMOS|8|1|主耶和华又指示我一件事，看哪，有一筐夏天的果子。
AMOS|8|2|他说：“ 阿摩司 ，你看见什么？”我说：“一筐夏天的果子。”耶和华对我说： “我子民 以色列 的结局 到了， 我必不再宽恕他们。
AMOS|8|3|那日，宫殿里的诗歌要变为哀号 ； 必有许多尸首抛在各处， 安静无声。” 这是主耶和华说的。
AMOS|8|4|你们这些践踏贫穷人、 使这地困苦人衰败的， 当听这话！
AMOS|8|5|你们说：“初一几时过去， 我们好卖粮； 安息日几时过去， 我们好摆开谷物； 我们要把伊法变小， 把舍客勒变大， 以诡诈的天平欺哄人，
AMOS|8|6|用银子买贫寒人， 以一双鞋换贫穷人， 把坏的谷物卖给人。”
AMOS|8|7|耶和华指着 雅各 的骄傲起誓说： “他们这一切的行为，我必永远不忘。
AMOS|8|8|地岂不因这事震动？ 其中的居民岂不悲哀吗？ 全地必如 尼罗河 涨起， 如 埃及 的 尼罗河 涌起退落。
AMOS|8|9|“到那日， 我要使太阳在正午落下， 使这地在白昼黑暗。” 这是主耶和华说的。
AMOS|8|10|“我要使你们的节期变为悲哀， 你们一切的歌曲变为哀歌； 我要使众人腰束麻布， 头上光秃； 我要使这悲哀如丧独子， 其结局如悲痛的日子。
AMOS|8|11|“看哪，日子将到， 我必命饥荒降在地上； 人饥饿非因无饼，干渴非因无水， 而是因不听耶和华的话。” 这是主耶和华说的。
AMOS|8|12|他们必飘流，从这海到那海， 从北边到东边，往来奔跑， 寻求耶和华的话， 却寻不着。
AMOS|8|13|“当那日，少年和美貌的少女 必因干渴而发昏。
AMOS|8|14|那些指着 撒玛利亚 的罪孽 起誓的，说： ‘ 但 哪，我们指着你那里的神明起誓’， 又说：‘我们指着通往 别是巴 的路起誓’， 这些人都必仆倒，永不再起。”
AMOS|9|1|我看见主站在祭坛旁，说： “你要击打柱顶，使门槛震动， 要剪除众人当中为首的， 他们中最后的 ，我必用刀杀戮； 无一人能逃避，无一人能逃脱。
AMOS|9|2|“虽然他们挖透阴间， 我的手必从那里拉出他们； 虽然他们爬到天上， 我必从那里拿下他们；
AMOS|9|3|虽然藏在 迦密山 顶， 我必在那里搜寻，擒拿他们； 虽然离开我眼前藏在海底， 我必在那里命令蛇咬他们；
AMOS|9|4|虽然被仇敌掳去， 我也必在那里命令刀剑杀戮他们； 我必定睛在他们身上， 降祸不降福。”
AMOS|9|5|万军的主耶和华触摸地，地就融化， 凡住在地上的都必悲哀； 全地必如 尼罗河 涨起， 如同 埃及 的 尼罗河 落下。
AMOS|9|6|那在天上建造楼阁、 在地上奠定穹苍、 召唤海水、 使其倾倒在地面上的， 耶和华是他的名。
AMOS|9|7|耶和华说：“ 以色列 人哪， 我岂不是看你们如 古实 人吗？ 我岂不是领 以色列 人出 埃及 地， 也领 非利士 人出 迦斐托 ， 领 亚兰 人出 吉珥 吗？
AMOS|9|8|看哪，主耶和华的眼目 察看这有罪的国度， 要把它从地面上灭绝， 却不将 雅各 家灭绝净尽。” 这是耶和华说的。
AMOS|9|9|“看哪，我发命令， 使 以色列 家在万国中飘流， 好像人用筛子筛谷， 连一粒也不落在地上。
AMOS|9|10|我子民中所有的罪人， 就是那些说 ‘灾祸必不靠近，必不追上我们’的， 都必死在刀下。”
AMOS|9|11|“在那日，我必重建 大卫 倒塌的帐幕， 修补其中的缺口； 我必建立那遭破坏的， 重新修造，如古时一般，
AMOS|9|12|使 以色列 人接管 以东 所剩余的 和所有称为我名下的国。 这是耶和华说的，他要行这事。
AMOS|9|13|“看哪，日子将到， 耕种的必接续收割的， 踹葡萄的必接续撒种的； 大山要滴下甜酒， 小山也被漫过。” 这是耶和华说的。
AMOS|9|14|“我要使 以色列 被掳的子民归回； 他们要重修荒废的城镇， 居住在其中； 栽植葡萄园，喝其中所出的酒， 修造果园，吃其中的果子。
AMOS|9|15|我要将他们栽植于本地， 他们必不再从我所赐给他们的地上被拔出。” 这是耶和华－你的上帝说的。
