2COR|1|1|Paul, an apostle of Christ Jesus by the will of God, and Timothy our brother, To the church of God in Corinth, together with all the saints throughout Achaia:
2COR|1|2|Grace and peace to you from God our Father and the Lord Jesus Christ.
2COR|1|3|Praise be to the God and Father of our Lord Jesus Christ, the Father of compassion and the God of all comfort,
2COR|1|4|who comforts us in all our troubles, so that we can comfort those in any trouble with the comfort we ourselves have received from God.
2COR|1|5|For just as the sufferings of Christ flow over into our lives, so also through Christ our comfort overflows.
2COR|1|6|If we are distressed, it is for your comfort and salvation; if we are comforted, it is for your comfort, which produces in you patient endurance of the same sufferings we suffer.
2COR|1|7|And our hope for you is firm, because we know that just as you share in our sufferings, so also you share in our comfort.
2COR|1|8|We do not want you to be uninformed, brothers, about the hardships we suffered in the province of Asia. We were under great pressure, far beyond our ability to endure, so that we despaired even of life.
2COR|1|9|Indeed, in our hearts we felt the sentence of death. But this happened that we might not rely on ourselves but on God, who raises the dead.
2COR|1|10|He has delivered us from such a deadly peril, and he will deliver us. On him we have set our hope that he will continue to deliver us,
2COR|1|11|as you help us by your prayers. Then many will give thanks on our behalf for the gracious favor granted us in answer to the prayers of many.
2COR|1|12|Now this is our boast: Our conscience testifies that we have conducted ourselves in the world, and especially in our relations with you, in the holiness and sincerity that are from God. We have done so not according to worldly wisdom but according to God's grace.
2COR|1|13|For we do not write you anything you cannot read or understand. And I hope that,
2COR|1|14|as you have understood us in part, you will come to understand fully that you can boast of us just as we will boast of you in the day of the Lord Jesus.
2COR|1|15|Because I was confident of this, I planned to visit you first so that you might benefit twice.
2COR|1|16|I planned to visit you on my way to Macedonia and to come back to you from Macedonia, and then to have you send me on my way to Judea.
2COR|1|17|When I planned this, did I do it lightly? Or do I make my plans in a worldly manner so that in the same breath I say, "Yes, yes" and "No, no"?
2COR|1|18|But as surely as God is faithful, our message to you is not "Yes" and "No."
2COR|1|19|For the Son of God, Jesus Christ, who was preached among you by me and Silas and Timothy, was not "Yes" and "No," but in him it has always been "Yes."
2COR|1|20|For no matter how many promises God has made, they are "Yes" in Christ. And so through him the "Amen" is spoken by us to the glory of God.
2COR|1|21|Now it is God who makes both us and you stand firm in Christ. He anointed us,
2COR|1|22|set his seal of ownership on us, and put his Spirit in our hearts as a deposit, guaranteeing what is to come.
2COR|1|23|I call God as my witness that it was in order to spare you that I did not return to Corinth.
2COR|1|24|Not that we lord it over your faith, but we work with you for your joy, because it is by faith you stand firm.
2COR|2|1|So I made up my mind that I would not make another painful visit to you.
2COR|2|2|For if I grieve you, who is left to make me glad but you whom I have grieved?
2COR|2|3|I wrote as I did so that when I came I should not be distressed by those who ought to make me rejoice. I had confidence in all of you, that you would all share my joy.
2COR|2|4|For I wrote you out of great distress and anguish of heart and with many tears, not to grieve you but to let you know the depth of my love for you.
2COR|2|5|If anyone has caused grief, he has not so much grieved me as he has grieved all of you, to some extent--not to put it too severely.
2COR|2|6|The punishment inflicted on him by the majority is sufficient for him.
2COR|2|7|Now instead, you ought to forgive and comfort him, so that he will not be overwhelmed by excessive sorrow.
2COR|2|8|I urge you, therefore, to reaffirm your love for him.
2COR|2|9|The reason I wrote you was to see if you would stand the test and be obedient in everything.
2COR|2|10|If you forgive anyone, I also forgive him. And what I have forgiven--if there was anything to forgive--I have forgiven in the sight of Christ for your sake,
2COR|2|11|in order that Satan might not outwit us. For we are not unaware of his schemes.
2COR|2|12|Now when I went to Troas to preach the gospel of Christ and found that the Lord had opened a door for me,
2COR|2|13|I still had no peace of mind, because I did not find my brother Titus there. So I said good-by to them and went on to Macedonia.
2COR|2|14|But thanks be to God, who always leads us in triumphal procession in Christ and through us spreads everywhere the fragrance of the knowledge of him.
2COR|2|15|For we are to God the aroma of Christ among those who are being saved and those who are perishing.
2COR|2|16|To the one we are the smell of death; to the other, the fragrance of life. And who is equal to such a task?
2COR|2|17|Unlike so many, we do not peddle the word of God for profit. On the contrary, in Christ we speak before God with sincerity, like men sent from God.
2COR|3|1|Are we beginning to commend ourselves again? Or do we need, like some people, letters of recommendation to you or from you?
2COR|3|2|You yourselves are our letter, written on our hearts, known and read by everybody.
2COR|3|3|You show that you are a letter from Christ, the result of our ministry, written not with ink but with the Spirit of the living God, not on tablets of stone but on tablets of human hearts.
2COR|3|4|Such confidence as this is ours through Christ before God.
2COR|3|5|Not that we are competent in ourselves to claim anything for ourselves, but our competence comes from God.
2COR|3|6|He has made us competent as ministers of a new covenant--not of the letter but of the Spirit; for the letter kills, but the Spirit gives life.
2COR|3|7|Now if the ministry that brought death, which was engraved in letters on stone, came with glory, so that the Israelites could not look steadily at the face of Moses because of its glory, fading though it was,
2COR|3|8|will not the ministry of the Spirit be even more glorious?
2COR|3|9|If the ministry that condemns men is glorious, how much more glorious is the ministry that brings righteousness!
2COR|3|10|For what was glorious has no glory now in comparison with the surpassing glory.
2COR|3|11|And if what was fading away came with glory, how much greater is the glory of that which lasts!
2COR|3|12|Therefore, since we have such a hope, we are very bold.
2COR|3|13|We are not like Moses, who would put a veil over his face to keep the Israelites from gazing at it while the radiance was fading away.
2COR|3|14|But their minds were made dull, for to this day the same veil remains when the old covenant is read. It has not been removed, because only in Christ is it taken away.
2COR|3|15|Even to this day when Moses is read, a veil covers their hearts.
2COR|3|16|But whenever anyone turns to the Lord, the veil is taken away.
2COR|3|17|Now the Lord is the Spirit, and where the Spirit of the Lord is, there is freedom.
2COR|3|18|And we, who with unveiled faces all reflect the Lord's glory, are being transformed into his likeness with ever-increasing glory, which comes from the Lord, who is the Spirit.
2COR|4|1|Therefore, since through God's mercy we have this ministry, we do not lose heart.
2COR|4|2|Rather, we have renounced secret and shameful ways; we do not use deception, nor do we distort the word of God. On the contrary, by setting forth the truth plainly we commend ourselves to every man's conscience in the sight of God.
2COR|4|3|And even if our gospel is veiled, it is veiled to those who are perishing.
2COR|4|4|The god of this age has blinded the minds of unbelievers, so that they cannot see the light of the gospel of the glory of Christ, who is the image of God.
2COR|4|5|For we do not preach ourselves, but Jesus Christ as Lord, and ourselves as your servants for Jesus' sake.
2COR|4|6|For God, who said, "Let light shine out of darkness," made his light shine in our hearts to give us the light of the knowledge of the glory of God in the face of Christ.
2COR|4|7|But we have this treasure in jars of clay to show that this all-surpassing power is from God and not from us.
2COR|4|8|We are hard pressed on every side, but not crushed; perplexed, but not in despair;
2COR|4|9|persecuted, but not abandoned; struck down, but not destroyed.
2COR|4|10|We always carry around in our body the death of Jesus, so that the life of Jesus may also be revealed in our body.
2COR|4|11|For we who are alive are always being given over to death for Jesus' sake, so that his life may be revealed in our mortal body.
2COR|4|12|So then, death is at work in us, but life is at work in you.
2COR|4|13|It is written: "I believed; therefore I have spoken." With that same spirit of faith we also believe and therefore speak,
2COR|4|14|because we know that the one who raised the Lord Jesus from the dead will also raise us with Jesus and present us with you in his presence.
2COR|4|15|All this is for your benefit, so that the grace that is reaching more and more people may cause thanksgiving to overflow to the glory of God.
2COR|4|16|Therefore we do not lose heart. Though outwardly we are wasting away, yet inwardly we are being renewed day by day.
2COR|4|17|For our light and momentary troubles are achieving for us an eternal glory that far outweighs them all.
2COR|4|18|So we fix our eyes not on what is seen, but on what is unseen. For what is seen is temporary, but what is unseen is eternal.
2COR|5|1|Now we know that if the earthly tent we live in is destroyed, we have a building from God, an eternal house in heaven, not built by human hands.
2COR|5|2|Meanwhile we groan, longing to be clothed with our heavenly dwelling,
2COR|5|3|because when we are clothed, we will not be found naked.
2COR|5|4|For while we are in this tent, we groan and are burdened, because we do not wish to be unclothed but to be clothed with our heavenly dwelling, so that what is mortal may be swallowed up by life.
2COR|5|5|Now it is God who has made us for this very purpose and has given us the Spirit as a deposit, guaranteeing what is to come.
2COR|5|6|Therefore we are always confident and know that as long as we are at home in the body we are away from the Lord.
2COR|5|7|We live by faith, not by sight.
2COR|5|8|We are confident, I say, and would prefer to be away from the body and at home with the Lord.
2COR|5|9|So we make it our goal to please him, whether we are at home in the body or away from it.
2COR|5|10|For we must all appear before the judgment seat of Christ, that each one may receive what is due him for the things done while in the body, whether good or bad.
2COR|5|11|Since, then, we know what it is to fear the Lord, we try to persuade men. What we are is plain to God, and I hope it is also plain to your conscience.
2COR|5|12|We are not trying to commend ourselves to you again, but are giving you an opportunity to take pride in us, so that you can answer those who take pride in what is seen rather than in what is in the heart.
2COR|5|13|If we are out of our mind, it is for the sake of God; if we are in our right mind, it is for you.
2COR|5|14|For Christ's love compels us, because we are convinced that one died for all, and therefore all died.
2COR|5|15|And he died for all, that those who live should no longer live for themselves but for him who died for them and was raised again.
2COR|5|16|So from now on we regard no one from a worldly point of view. Though we once regarded Christ in this way, we do so no longer.
2COR|5|17|Therefore, if anyone is in Christ, he is a new creation; the old has gone, the new has come!
2COR|5|18|All this is from God, who reconciled us to himself through Christ and gave us the ministry of reconciliation:
2COR|5|19|that God was reconciling the world to himself in Christ, not counting men's sins against them. And he has committed to us the message of reconciliation.
2COR|5|20|We are therefore Christ's ambassadors, as though God were making his appeal through us. We implore you on Christ's behalf: Be reconciled to God.
2COR|5|21|God made him who had no sin to be sin for us, so that in him we might become the righteousness of God.
2COR|6|1|As God's fellow workers we urge you not to receive God's grace in vain.
2COR|6|2|For he says, "In the time of my favor I heard you, and in the day of salvation I helped you." I tell you, now is the time of God's favor, now is the day of salvation.
2COR|6|3|We put no stumbling block in anyone's path, so that our ministry will not be discredited.
2COR|6|4|Rather, as servants of God we commend ourselves in every way: in great endurance; in troubles, hardships and distresses;
2COR|6|5|in beatings, imprisonments and riots; in hard work, sleepless nights and hunger;
2COR|6|6|in purity, understanding, patience and kindness; in the Holy Spirit and in sincere love;
2COR|6|7|in truthful speech and in the power of God; with weapons of righteousness in the right hand and in the left;
2COR|6|8|through glory and dishonor, bad report and good report; genuine, yet regarded as impostors;
2COR|6|9|known, yet regarded as unknown; dying, and yet we live on; beaten, and yet not killed;
2COR|6|10|sorrowful, yet always rejoicing; poor, yet making many rich; having nothing, and yet possessing everything.
2COR|6|11|We have spoken freely to you, Corinthians, and opened wide our hearts to you.
2COR|6|12|We are not withholding our affection from you, but you are withholding yours from us.
2COR|6|13|As a fair exchange--I speak as to my children--open wide your hearts also.
2COR|6|14|Do not be yoked together with unbelievers. For what do righteousness and wickedness have in common? Or what fellowship can light have with darkness?
2COR|6|15|What harmony is there between Christ and Belial? What does a believer have in common with an unbeliever?
2COR|6|16|What agreement is there between the temple of God and idols? For we are the temple of the living God. As God has said: "I will live with them and walk among them, and I will be their God, and they will be my people."
2COR|6|17|"Therefore come out from them and be separate, says the Lord. Touch no unclean thing, and I will receive you."
2COR|6|18|"I will be a Father to you, and you will be my sons and daughters, says the Lord Almighty."
2COR|7|1|Since we have these promises, dear friends, let us purify ourselves from everything that contaminates body and spirit, perfecting holiness out of reverence for God.
2COR|7|2|Make room for us in your hearts. We have wronged no one, we have corrupted no one, we have exploited no one.
2COR|7|3|I do not say this to condemn you; I have said before that you have such a place in our hearts that we would live or die with you.
2COR|7|4|I have great confidence in you; I take great pride in you. I am greatly encouraged; in all our troubles my joy knows no bounds.
2COR|7|5|For when we came into Macedonia, this body of ours had no rest, but we were harassed at every turn--conflicts on the outside, fears within.
2COR|7|6|But God, who comforts the downcast, comforted us by the coming of Titus,
2COR|7|7|and not only by his coming but also by the comfort you had given him. He told us about your longing for me, your deep sorrow, your ardent concern for me, so that my joy was greater than ever.
2COR|7|8|Even if I caused you sorrow by my letter, I do not regret it. Though I did regret it--I see that my letter hurt you, but only for a little while--
2COR|7|9|yet now I am happy, not because you were made sorry, but because your sorrow led you to repentance. For you became sorrowful as God intended and so were not harmed in any way by us.
2COR|7|10|Godly sorrow brings repentance that leads to salvation and leaves no regret, but worldly sorrow brings death.
2COR|7|11|See what this godly sorrow has produced in you: what earnestness, what eagerness to clear yourselves, what indignation, what alarm, what longing, what concern, what readiness to see justice done. At every point you have proved yourselves to be innocent in this matter.
2COR|7|12|So even though I wrote to you, it was not on account of the one who did the wrong or of the injured party, but rather that before God you could see for yourselves how devoted to us you are.
2COR|7|13|By all this we are encouraged.
2COR|7|14|In addition to our own encouragement, we were especially delighted to see how happy Titus was, because his spirit has been refreshed by all of you. I had boasted to him about you, and you have not embarrassed me. But just as everything we said to you was true, so our boasting about you to Titus has proved to be true as well.
2COR|7|15|And his affection for you is all the greater when he remembers that you were all obedient, receiving him with fear and trembling.
2COR|7|16|I am glad I can have complete confidence in you.
2COR|8|1|And now, brothers, we want you to know about the grace that God has given the Macedonian churches.
2COR|8|2|Out of the most severe trial, their overflowing joy and their extreme poverty welled up in rich generosity.
2COR|8|3|For I testify that they gave as much as they were able, and even beyond their ability. Entirely on their own,
2COR|8|4|they urgently pleaded with us for the privilege of sharing in this service to the saints.
2COR|8|5|And they did not do as we expected, but they gave themselves first to the Lord and then to us in keeping with God's will.
2COR|8|6|So we urged Titus, since he had earlier made a beginning, to bring also to completion this act of grace on your part.
2COR|8|7|But just as you excel in everything--in faith, in speech, in knowledge, in complete earnestness and in your love for us--see that you also excel in this grace of giving.
2COR|8|8|I am not commanding you, but I want to test the sincerity of your love by comparing it with the earnestness of others.
2COR|8|9|For you know the grace of our Lord Jesus Christ, that though he was rich, yet for your sakes he became poor, so that you through his poverty might become rich.
2COR|8|10|And here is my advice about what is best for you in this matter: Last year you were the first not only to give but also to have the desire to do so.
2COR|8|11|Now finish the work, so that your eager willingness to do it may be matched by your completion of it, according to your means.
2COR|8|12|For if the willingness is there, the gift is acceptable according to what one has, not according to what he does not have.
2COR|8|13|Our desire is not that others might be relieved while you are hard pressed, but that there might be equality.
2COR|8|14|At the present time your plenty will supply what they need, so that in turn their plenty will supply what you need. Then there will be equality,
2COR|8|15|as it is written: "He who gathered much did not have too much, and he who gathered little did not have too little."
2COR|8|16|I thank God, who put into the heart of Titus the same concern I have for you.
2COR|8|17|For Titus not only welcomed our appeal, but he is coming to you with much enthusiasm and on his own initiative.
2COR|8|18|And we are sending along with him the brother who is praised by all the churches for his service to the gospel.
2COR|8|19|What is more, he was chosen by the churches to accompany us as we carry the offering, which we administer in order to honor the Lord himself and to show our eagerness to help.
2COR|8|20|We want to avoid any criticism of the way we administer this liberal gift.
2COR|8|21|For we are taking pains to do what is right, not only in the eyes of the Lord but also in the eyes of men.
2COR|8|22|In addition, we are sending with them our brother who has often proved to us in many ways that he is zealous, and now even more so because of his great confidence in you.
2COR|8|23|As for Titus, he is my partner and fellow worker among you; as for our brothers, they are representatives of the churches and an honor to Christ.
2COR|8|24|Therefore show these men the proof of your love and the reason for our pride in you, so that the churches can see it.
2COR|9|1|There is no need for me to write to you about this service to the saints.
2COR|9|2|For I know your eagerness to help, and I have been boasting about it to the Macedonians, telling them that since last year you in Achaia were ready to give; and your enthusiasm has stirred most of them to action.
2COR|9|3|But I am sending the brothers in order that our boasting about you in this matter should not prove hollow, but that you may be ready, as I said you would be.
2COR|9|4|For if any Macedonians come with me and find you unprepared, we--not to say anything about you--would be ashamed of having been so confident.
2COR|9|5|So I thought it necessary to urge the brothers to visit you in advance and finish the arrangements for the generous gift you had promised. Then it will be ready as a generous gift, not as one grudgingly given.
2COR|9|6|Remember this: Whoever sows sparingly will also reap sparingly, and whoever sows generously will also reap generously.
2COR|9|7|Each man should give what he has decided in his heart to give, not reluctantly or under compulsion, for God loves a cheerful giver.
2COR|9|8|And God is able to make all grace abound to you, so that in all things at all times, having all that you need, you will abound in every good work.
2COR|9|9|As it is written: "He has scattered abroad his gifts to the poor; his righteousness endures forever."
2COR|9|10|Now he who supplies seed to the sower and bread for food will also supply and increase your store of seed and will enlarge the harvest of your righteousness.
2COR|9|11|You will be made rich in every way so that you can be generous on every occasion, and through us your generosity will result in thanksgiving to God.
2COR|9|12|This service that you perform is not only supplying the needs of God's people but is also overflowing in many expressions of thanks to God.
2COR|9|13|Because of the service by which you have proved yourselves, men will praise God for the obedience that accompanies your confession of the gospel of Christ, and for your generosity in sharing with them and with everyone else.
2COR|9|14|And in their prayers for you their hearts will go out to you, because of the surpassing grace God has given you.
2COR|9|15|Thanks be to God for his indescribable gift!
2COR|10|1|By the meekness and gentleness of Christ, I appeal to you--I, Paul, who am "timid" when face to face with you, but "bold" when away!
2COR|10|2|I beg you that when I come I may not have to be as bold as I expect to be toward some people who think that we live by the standards of this world.
2COR|10|3|For though we live in the world, we do not wage war as the world does.
2COR|10|4|The weapons we fight with are not the weapons of the world. On the contrary, they have divine power to demolish strongholds.
2COR|10|5|We demolish arguments and every pretension that sets itself up against the knowledge of God, and we take captive every thought to make it obedient to Christ.
2COR|10|6|And we will be ready to punish every act of disobedience, once your obedience is complete.
2COR|10|7|You are looking only on the surface of things. If anyone is confident that he belongs to Christ, he should consider again that we belong to Christ just as much as he.
2COR|10|8|For even if I boast somewhat freely about the authority the Lord gave us for building you up rather than pulling you down, I will not be ashamed of it.
2COR|10|9|I do not want to seem to be trying to frighten you with my letters.
2COR|10|10|For some say, "His letters are weighty and forceful, but in person he is unimpressive and his speaking amounts to nothing."
2COR|10|11|Such people should realize that what we are in our letters when we are absent, we will be in our actions when we are present.
2COR|10|12|We do not dare to classify or compare ourselves with some who commend themselves. When they measure themselves by themselves and compare themselves with themselves, they are not wise.
2COR|10|13|We, however, will not boast beyond proper limits, but will confine our boasting to the field God has assigned to us, a field that reaches even to you.
2COR|10|14|We are not going too far in our boasting, as would be the case if we had not come to you, for we did get as far as you with the gospel of Christ.
2COR|10|15|Neither do we go beyond our limits by boasting of work done by others. Our hope is that, as your faith continues to grow, our area of activity among you will greatly expand,
2COR|10|16|so that we can preach the gospel in the regions beyond you. For we do not want to boast about work already done in another man's territory.
2COR|10|17|But, "Let him who boasts boast in the Lord."
2COR|10|18|For it is not the one who commends himself who is approved, but the one whom the Lord commends.
2COR|11|1|I hope you will put up with a little of my foolishness; but you are already doing that.
2COR|11|2|I am jealous for you with a godly jealousy. I promised you to one husband, to Christ, so that I might present you as a pure virgin to him.
2COR|11|3|But I am afraid that just as Eve was deceived by the serpent's cunning, your minds may somehow be led astray from your sincere and pure devotion to Christ.
2COR|11|4|For if someone comes to you and preaches a Jesus other than the Jesus we preached, or if you receive a different spirit from the one you received, or a different gospel from the one you accepted, you put up with it easily enough.
2COR|11|5|But I do not think I am in the least inferior to those "super-apostles."
2COR|11|6|I may not be a trained speaker, but I do have knowledge. We have made this perfectly clear to you in every way.
2COR|11|7|Was it a sin for me to lower myself in order to elevate you by preaching the gospel of God to you free of charge?
2COR|11|8|I robbed other churches by receiving support from them so as to serve you.
2COR|11|9|And when I was with you and needed something, I was not a burden to anyone, for the brothers who came from Macedonia supplied what I needed. I have kept myself from being a burden to you in any way, and will continue to do so.
2COR|11|10|As surely as the truth of Christ is in me, nobody in the regions of Achaia will stop this boasting of mine.
2COR|11|11|Why? Because I do not love you? God knows I do!
2COR|11|12|And I will keep on doing what I am doing in order to cut the ground from under those who want an opportunity to be considered equal with us in the things they boast about.
2COR|11|13|For such men are false apostles, deceitful workmen, masquerading as apostles of Christ.
2COR|11|14|And no wonder, for Satan himself masquerades as an angel of light.
2COR|11|15|It is not surprising, then, if his servants masquerade as servants of righteousness. Their end will be what their actions deserve.
2COR|11|16|I repeat: Let no one take me for a fool. But if you do, then receive me just as you would a fool, so that I may do a little boasting.
2COR|11|17|In this self-confident boasting I am not talking as the Lord would, but as a fool.
2COR|11|18|Since many are boasting in the way the world does, I too will boast.
2COR|11|19|You gladly put up with fools since you are so wise!
2COR|11|20|In fact, you even put up with anyone who enslaves you or exploits you or takes advantage of you or pushes himself forward or slaps you in the face.
2COR|11|21|To my shame I admit that we were too weak for that!
2COR|11|22|What anyone else dares to boast about--I am speaking as a fool--I also dare to boast about. Are they Hebrews? So am I. Are they Israelites? So am I. Are they Abraham's descendants? So am I.
2COR|11|23|Are they servants of Christ? (I am out of my mind to talk like this.) I am more. I have worked much harder, been in prison more frequently, been flogged more severely, and been exposed to death again and again.
2COR|11|24|Five times I received from the Jews the forty lashes minus one.
2COR|11|25|Three times I was beaten with rods, once I was stoned, three times I was shipwrecked, I spent a night and a day in the open sea,
2COR|11|26|I have been constantly on the move. I have been in danger from rivers, in danger from bandits, in danger from my own countrymen, in danger from Gentiles; in danger in the city, in danger in the country, in danger at sea; and in danger from false brothers.
2COR|11|27|I have labored and toiled and have often gone without sleep; I have known hunger and thirst and have often gone without food; I have been cold and naked.
2COR|11|28|Besides everything else, I face daily the pressure of my concern for all the churches.
2COR|11|29|Who is weak, and I do not feel weak? Who is led into sin, and I do not inwardly burn?
2COR|11|30|If I must boast, I will boast of the things that show my weakness.
2COR|11|31|The God and Father of the Lord Jesus, who is to be praised forever, knows that I am not lying.
2COR|11|32|In Damascus the governor under King Aretas had the city of the Damascenes guarded in order to arrest me.
2COR|11|33|But I was lowered in a basket from a window in the wall and slipped through his hands.
2COR|12|1|I must go on boasting. Although there is nothing to be gained, I will go on to visions and revelations from the Lord.
2COR|12|2|I know a man in Christ who fourteen years ago was caught up to the third heaven. Whether it was in the body or out of the body I do not know--God knows.
2COR|12|3|And I know that this man--whether in the body or apart from the body I do not know, but God knows--
2COR|12|4|was caught up to paradise. He heard inexpressible things, things that man is not permitted to tell.
2COR|12|5|I will boast about a man like that, but I will not boast about myself, except about my weaknesses.
2COR|12|6|Even if I should choose to boast, I would not be a fool, because I would be speaking the truth. But I refrain, so no one will think more of me than is warranted by what I do or say.
2COR|12|7|To keep me from becoming conceited because of these surpassingly great revelations, there was given me a thorn in my flesh, a messenger of Satan, to torment me.
2COR|12|8|Three times I pleaded with the Lord to take it away from me.
2COR|12|9|But he said to me, "My grace is sufficient for you, for my power is made perfect in weakness." Therefore I will boast all the more gladly about my weaknesses, so that Christ's power may rest on me.
2COR|12|10|That is why, for Christ's sake, I delight in weaknesses, in insults, in hardships, in persecutions, in difficulties. For when I am weak, then I am strong.
2COR|12|11|I have made a fool of myself, but you drove me to it. I ought to have been commended by you, for I am not in the least inferior to the "super-apostles," even though I am nothing.
2COR|12|12|The things that mark an apostle--signs, wonders and miracles--were done among you with great perseverance.
2COR|12|13|How were you inferior to the other churches, except that I was never a burden to you? Forgive me this wrong!
2COR|12|14|Now I am ready to visit you for the third time, and I will not be a burden to you, because what I want is not your possessions but you. After all, children should not have to save up for their parents, but parents for their children.
2COR|12|15|So I will very gladly spend for you everything I have and expend myself as well. If I love you more, will you love me less?
2COR|12|16|Be that as it may, I have not been a burden to you. Yet, crafty fellow that I am, I caught you by trickery!
2COR|12|17|Did I exploit you through any of the men I sent you?
2COR|12|18|I urged Titus to go to you and I sent our brother with him. Titus did not exploit you, did he? Did we not act in the same spirit and follow the same course?
2COR|12|19|Have you been thinking all along that we have been defending ourselves to you? We have been speaking in the sight of God as those in Christ; and everything we do, dear friends, is for your strengthening.
2COR|12|20|For I am afraid that when I come I may not find you as I want you to be, and you may not find me as you want me to be. I fear that there may be quarreling, jealousy, outbursts of anger, factions, slander, gossip, arrogance and disorder.
2COR|12|21|I am afraid that when I come again my God will humble me before you, and I will be grieved over many who have sinned earlier and have not repented of the impurity, sexual sin and debauchery in which they have indulged.
2COR|13|1|This will be my third visit to you. "Every matter must be established by the testimony of two or three witnesses."
2COR|13|2|I already gave you a warning when I was with you the second time. I now repeat it while absent: On my return I will not spare those who sinned earlier or any of the others,
2COR|13|3|since you are demanding proof that Christ is speaking through me. He is not weak in dealing with you, but is powerful among you.
2COR|13|4|For to be sure, he was crucified in weakness, yet he lives by God's power. Likewise, we are weak in him, yet by God's power we will live with him to serve you.
2COR|13|5|Examine yourselves to see whether you are in the faith; test yourselves. Do you not realize that Christ Jesus is in you--unless, of course, you fail the test?
2COR|13|6|And I trust that you will discover that we have not failed the test.
2COR|13|7|Now we pray to God that you will not do anything wrong. Not that people will see that we have stood the test but that you will do what is right even though we may seem to have failed.
2COR|13|8|For we cannot do anything against the truth, but only for the truth.
2COR|13|9|We are glad whenever we are weak but you are strong; and our prayer is for your perfection.
2COR|13|10|This is why I write these things when I am absent, that when I come I may not have to be harsh in my use of authority--the authority the Lord gave me for building you up, not for tearing you down.
2COR|13|11|Finally, brothers, good-by. Aim for perfection, listen to my appeal, be of one mind, live in peace. And the God of love and peace will be with you.
2COR|13|12|Greet one another with a holy kiss.
2COR|13|13|All the saints send their greetings.
2COR|13|14|May the grace of the Lord Jesus Christ, and the love of God, and the fellowship of the Holy Spirit be with you all.
