ECCL|1|1|Verba Ecclesiastes filii David regis Ierusalem."
ECCL|1|2|" Vanitas vanitatum,dixit Ecclesiastes,vanitas vanitatum et omnia vanitas ".
ECCL|1|3|Quid lucri est hominide universo labore suo, quo laborat sub sole?
ECCL|1|4|Generatio praeterit, et generatio advenit,terra autem in aeternum stat.
ECCL|1|5|Oritur sol, et occidit solet ad locum suum anhelat ibique renascitur.
ECCL|1|6|Gyrat per meridiem et flectitur ad aquilonem,lustrans universa in circuitu pergit spirituset in circulos suos revertitur.
ECCL|1|7|Omnia flumina pergunt ad mare, et mare non redundat;ad locum, unde exeunt, flumina illuc revertuntur in cursu suo.
ECCL|1|8|Cunctae res difficiles;non potest eas homo explicare sermone.Non saturatur oculus visu,nec auris auditu impletur.
ECCL|1|9|Quod fuit,ipsum est, quod futurum est.Quod factum est,ipsum est, quod faciendum est:
ECCL|1|10|nihil sub sole novum.Si de quadam re dicitur: " Ecce hoc novum est ",iam enim praecessit in saeculis, quae fuerunt ante nos.
ECCL|1|11|Non est priorum memoria,sed nec eorum quidem, qui postea futuri sunt,erit recordatio apud eos,qui futuri sunt in novissimo.
ECCL|1|12|Ego Ecclesiastes fui rex Israel in Ierusalem
ECCL|1|13|et proposui in animo meo quaerere et investigare sapienter de omnibus, quae fiunt sub sole. Hanc occupationem pessimam dedit Deus filiis hominum, ut occuparentur in ea.
ECCL|1|14|Vidi cuncta, quae fiunt sub sole; et ecce universa vanitas et afflictio spiritus.
ECCL|1|15|Quod est curvum, rectum fieri non potest;et, quod deficiens est, numerari non potest.
ECCL|1|16|Locutus sum ego in corde meo dicens: " Ecce ego magnificavi et apposui sapientiam super omnes, qui fuerunt ante me in Ierusalem; et mens mea contemplata est multam sapientiam et scientiam ".
ECCL|1|17|Dedique cor meum, ut scirem sapientiam et scientiam, insipientiam et stultitiam. Et agnovi quod in his quoque esset afflictio spiritus, eo quod
ECCL|1|18|in multa sapientia multus sit maeror;et, qui addit scientiam, addit et laborem.
ECCL|2|1|Dixi ego in corde meo: " Veni, tentabo te gaudio: fruere bo nis "; et ecce hoc quoque vanitas.
ECCL|2|2|De risu dixi: " Insania "et de gaudio: " Quid prodest? ".
ECCL|2|3|Tractavi in corde meo detinere in vino carnem meam, cum cor meum duceretur in sapientia, et amplecti stultitiam, donec viderem quid esset utile filiis hominum, ut faciant sub sole paucis diebus vitae suae.
ECCL|2|4|Magnificavi opera mea: aedificavi mihi domos et plantavi vineas,
ECCL|2|5|feci hortos et pomaria et consevi ea arboribus cuncti generis fructuum
ECCL|2|6|et exstruxi mihi piscinas aquarum, ut irrigarem silvam lignorum germinantium.
ECCL|2|7|Possedi servos et ancillas et habui multam familiam, habui armenta quoque et magnos ovium greges ultra omnes, qui fuerunt ante me in Ierusalem.
ECCL|2|8|Coacervavi mihi etiam argentum et aurum et substantias regum ac provinciarum, feci mihi cantores et cantatrices et delicias filiorum hominum, scyphos et urceos in ministerio ad vina fundenda
ECCL|2|9|et crevi, supergressus sum omnes, qui ante me fuerunt in Ierusalem; sapientia quoque mea perseveravit mecum.
ECCL|2|10|Et omnia, quae desideraverunt oculi mei, non negavi eis nec prohibui cor meum ab omni voluptate, et oblectatum est ex omnibus laboribus, et hanc ratus sum partem meam ab omnibus aerumnis meis.
ECCL|2|11|Cumque me convertissem ad universa opera, quae fecerant manus meae, et ad labores, in quibus sudaveram, et ecce in omnibus vanitas et afflictio spiritus, et nihil lucri esse sub sole.
ECCL|2|12|Verti me ad contemplandam sapientiam et insipientiam et stultitiam: " Quid faciet, inquam, homo, qui veniet post regem? Id quod antea fecerunt.
ECCL|2|13|Et vidi quod tantum praecederet sapientia stultitiam, quantum lux praecedit tenebras.
ECCL|2|14|" Sapientis oculi in capite eius,stultus in tenebris ambulat ";et didici quod unus utriusqueesset interitus.
ECCL|2|15|Et dixi in corde meo: " Si unus et stulti et meus occasus erit, quid mihi prodest quod maiorem sapientiae dedi operam? ". Locutusque cum mente mea, animadverti quod hoc quoque esset vanitas.
ECCL|2|16|Non enim erit memoria sapientis similiter ut stulti in perpetuum; siquidem futura tempora oblivione cuncta pariter operient: moritur doctus similiter ut indoctus.
ECCL|2|17|Et idcirco taeduit me vitae meae, quia malum mihi est, quod sub sole fit; cuncta enim vanitas et afflictio spiritus.
ECCL|2|18|Rursus detestatus sum omnem laborem meum, quo sub sole laboravi, quem relicturus sum homini, qui erit post me;
ECCL|2|19|et quis scit utrum sapiens an stultus futurus sit? Et dominabitur in laboribus meis, quibus desudavi et sollicitus fui sub sole. Hoc quoque vanitas.
ECCL|2|20|Verti me exasperans cor meum de omni labore, quo laboravi sub sole.
ECCL|2|21|Nam est qui laborat in sapientia et doctrina et sollicitudine, et homini, qui non laboraverit, dabit portionem suam; et hoc ergo vanitas et magnum malum.
ECCL|2|22|Quid enim proderit homini de universo labore suo et afflictione cordis, qua sub sole laboravit?
ECCL|2|23|Cuncti dies eius dolores sunt, et aerumnae occupatio eius, nec per noctem cor eius requiescit; et hoc quoque vanitas est.
ECCL|2|24|Nihil melius est homini quam comedere et bibere et ostendere animae suae bona de laboribus suis. Et hoc vidi de manu Dei esse.
ECCL|2|25|Quis enim comedet et deliciis affluet sine eo?
ECCL|2|26|Quia homini bono in conspectu suo dedit sapientiam et scientiam et laetitiam; peccatori autem dedit afflictionem colligendi et congregandi, ut tradat ei, qui placuit Deo; sed et hoc vanitas est et afflictio spiritus.
ECCL|3|1|Omnia tempus habent,et momentum suum cuique negotio sub caelo:
ECCL|3|2|tempus nascendi et tempus moriendi,tempus plantandi et tempus evellendi quod plantatum est,
ECCL|3|3|tempus occidendi et tempus sanandi,tempus destruendi et tempus aedificandi,
ECCL|3|4|tempus flendi et tempus ridendi,tempus plangendi et tempus saltandi,
ECCL|3|5|tempus spargendi lapides et tempus eos colligendi,tempus amplexandi et tempus longe fieri ab amplexibus,
ECCL|3|6|tempus quaerendi et tempus perdendi,tempus custodiendi et tempus abiciendi,
ECCL|3|7|tempus scindendi et tempus consuendi,tempus tacendi et tempus loquendi,
ECCL|3|8|tempus dilectionis et tempus odii,tempus belli et tempus pacis.
ECCL|3|9|Quid lucri habet, qui operatur, de labore suo?
ECCL|3|10|Vidi occupationem, quam dedit Deus filiis hominum, ut occuparentur in ea.
ECCL|3|11|Cuncta fecit bona in tempore suo; et mundum tradidit cordi eorum, et non inveniet homo opus, quod operatus est Deus ab initio usque ad finem.
ECCL|3|12|Cognovi quod nihil boni esset in eis nisi laetari et facere bene in vita sua.
ECCL|3|13|Omnis enim homo, qui comedit et bibit et videt bonum de labore suo, hoc donum Dei est.
ECCL|3|14|Didici quod omnia opera, quae fecit Deus, perseverent in perpetuum; non possumus eis quidquam addere nec auferre, quae fecit Deus, ut timeatur.
ECCL|3|15|Quod iam fuit, ipsum est; et, quod futurum est, iam fuit; et Deus requirit, quod abiit.
ECCL|3|16|Et adhuc vidi sub sole: in loco iudicii ibi impietas, et in loco iustitiae ibi iniquitas;
ECCL|3|17|et dixi in corde meo: " Iustum et impium iudicabit Deus, quia tempus omni rei et omnibus occasio ".
ECCL|3|18|Dixi in corde meo de filiis hominum, ut probaret eos Deus et ostenderet eos in semetipsis similes esse bestiis.
ECCL|3|19|Quoniam sors filiorum hominis et iumentorum una est atque eadem: sicut moritur homo, sic et illa moriuntur; et idem spiritus omnibus: nihil habet homo iumento amplius, quia omnia vanitas.
ECCL|3|20|Et omnia pergunt ad unum locum:de terra facta sunt omnia,et in terram omnia pariter revertuntur.
ECCL|3|21|Quis novit, si spiritus filiorum hominis ascendat sursum, et si spiritus iumentorum descendat deorsum in terram?
ECCL|3|22|Et deprehendi nihil esse melius quam laetari hominem in opere suo; nam haec est pars illius. Quis enim eum adducet, ut post se futura cognoscat?
ECCL|4|1|Verti me ad alia et vidi calumnias, quae sub sole geruntur, et ecce lacrimae oppressorum, et nemo consolator; et ex parte opprimentium violentia, et nemo consolator.
ECCL|4|2|Et laudavi magis mortuos, qui iam defuncti sunt, quam viventes, qui adhuc vitam agunt,
ECCL|4|3|et feliciorem utroque iudicavi, qui necdum natus est nec vidit opera mala, quae sub sole fiunt.
ECCL|4|4|Rursum contemplatus sum omnes labores et omnem successum operis, et hoc esse zelum in proximum suum. Et in hoc ergo vanitas et afflictio spiritus.
ECCL|4|5|Stultus complicat manus suaset comedit carnes suas.
ECCL|4|6|Melior est pugillus cum requiequam plena utraque manus cum labore et afflictione spiritus.
ECCL|4|7|Iterum repperi et aliam vanitatem sub sole:
ECCL|4|8|unus est et secundum non habet, non filium, non fratrem, et tamen laborare non cessat, nec satiantur oculi eius divitiis, nec recogitat dicens: " Cui laboro et fraudo animam meam bonis?". In hoc quoque vanitas est et occupatio pessima.
ECCL|4|9|Melius est duos esse simul quam unum: habent enim emolumentum in labore suo,
ECCL|4|10|quia si unus ceciderit, ab altero fulcietur. Vae soli! Cum ceciderit, non habet sublevantem se.
ECCL|4|11|Insuper, si dormierint duo, fovebuntur mutuo; unus quomodo calefiet?
ECCL|4|12|Et, si quispiam praevaluerit contra unum, duo resistent ei. Et fu niculus triplex non cito rumpitur.
ECCL|4|13|Melior est puer pauper et sapiensrege sene et stulto,qui iam nescit erudiri.
ECCL|4|14|Ille enim de domo carceris exivit, ut regnaret, etiamsi in regno istius natus sit pauper.
ECCL|4|15|Vidi cunctos viventes, qui ambulant sub sole, cum adulescente illo secundo, qui consurgebat pro eo.
ECCL|4|16|Infinitus numerus erat populi, omnium, quos ipse praecedebat; sed qui postea futuri sunt, non laetabuntur in eo. Et hoc vanitas et afflictio spiritus.
ECCL|4|17|Custodi pedem tuum ingrediens domum Dei, nam accedere, ut audias, melius est quam cum stulti offerunt victimas: multo enim melior est oboedientia quam stultorum victimae, qui nesciunt se malum facere.
ECCL|5|1|Ne temere quid loquaris, neque cor tuum sit velox ad proferen dum sermonem coram Deo; Deus enim in caelo, et tu super terram: idcirco sint pauci sermones tui.
ECCL|5|2|Multas curas sequuntur somnia,et in multis sermonibus invenietur stultitia.
ECCL|5|3|Si quid vovisti Deo, ne moreris reddere: displicet enim ei stulta promissio; sed, quodcumque voveris, redde.
ECCL|5|4|Multoque melius est non vovere, quam post votum promissa non reddere.
ECCL|5|5|Ne dederis os tuum, ut peccare faciat carnem tuam, neque dicas coram angelo: " Error fuit "; ne forte iratus Deus contra sermones tuos dissipet opera manuum tuarum.
ECCL|5|6|Ubi multa sunt somnia, plurimae sunt vanitates et sermones innumeri; tu vero Deum time.
ECCL|5|7|Si videris calumnias egenorum et subreptionem iudicii et iustitiae in provincia, non mireris super hoc negotio, quia excelso excelsior vigilat, et super hos quoque eminentiores sunt alii;
ECCL|5|8|et terrae lucrum in omnibus est rex, cuius agri culti sunt.
ECCL|5|9|Qui diligit pecuniam, pecunia non implebitur; et, qui amat divitias, fructum non capiet ex eis; et hoc ergo vanitas.
ECCL|5|10|Ubi multae sunt opes, multi et qui comedunt eas; et quid prodest possessori, nisi quod cernit divitias oculis suis?
ECCL|5|11|Dulcis est somnus operanti,sive parum sive multum comedat;saturitas autem divitisnon sinit eum dormire.
ECCL|5|12|Est et infirmitas pessima, quam vidi sub sole: divitiae conservatae in malum domini sui.
ECCL|5|13|Perierunt enim in negotio pessimo; si generavit filium, in summa egestate erit.
ECCL|5|14|Sicut egressus est de utero matris suae, nudus iterum abibit, sicut venit, et nihil auferet secum de labore suo, quod tollat in manu sua.
ECCL|5|15|Miserabilis prorsus infirmitas: quomodo venit, sic revertetur. Quid ergo prodest ei quod laboravit in ventum?
ECCL|5|16|Cunctis enim diebus vitae suae comedit in tenebris et in curis multis et in aerumna atque tristitia.
ECCL|5|17|Ecce quod ego vidi bonum, quod pulchrum, ut comedat quis et bibat et fruatur laetitia ex labore suo, quo laboravit ipse sub sole, numero dierum vitae suae, quos dedit ei Deus; haec enim est pars illius.
ECCL|5|18|Et quidem omni homini, cui dedit Deus divitias atque substantiam, potestatemque ei tribuit, ut comedat ex eis et tollat partem suam et laetetur de labore suo: hoc est donum Dei.
ECCL|5|19|Non enim satis recordabitur dierum vitae suae, eo quod Deus occupet deliciis cor eius.
ECCL|6|1|Est et aliud malum, quod vidi sub sole, et quidem grave apud homines:
ECCL|6|2|vir, cui dedit Deus divitias et substantiam et honorem, et nihil deest animae suae ex omnibus, quae desiderat; nec tribuit ei potestatem Deus, ut comedat ex eo, sed homo extraneus vorabit illud: hoc vanitas et miseria mala est.
ECCL|6|3|Si genuerit quispiam centum liberos et vixerit multos annos et plures dies aetatis habuerit, et anima illius non sit satiata bonis substantiae suae, immo et sepultura careat, de hoc ego pronuntio quod melior illo sit abortivus.
ECCL|6|4|Frustra enim venit et pergit ad tenebras, et in tenebris abscondetur nomen eius.
ECCL|6|5|Etsi non vidit solem neque cognovit, maior est requies isti quam illi.
ECCL|6|6|Etiamsi duobus milibus annis vixerit et non fuerit perfruitus bonis, nonne ad unum locum properant omnes?
ECCL|6|7|" Omnis labor hominis est ad os eius,sed anima eius non implebitur ".
ECCL|6|8|Quid habet amplius sapiens prae stulto? Et quid pauper, qui sciat ambulare coram vivis?
ECCL|6|9|" Melior est oculorum visio quam vana persequi desideria "; sed et hoc vanitas est et afflictio spiritus.
ECCL|6|10|Quidquid est, iam vocatum est nomen eius; et scitur quod homo sit et non possit contra fortiorem se in iudicio contendere.
ECCL|6|11|Ubi verba sunt plurima, multiplicant vanitatem; quid lucri habet homo?
ECCL|6|12|Quoniam quis scit quid homini bonum sit in vita, in paucis diebus vanitatis suae, quos peragit velut umbra? Aut quis ei poterit indicare quid post eum futurum sub sole sit?
ECCL|7|1|Melius est nomen bonum quam unguenta pretiosa,et dies mortis die nativitatis.
ECCL|7|2|Melius est ire ad domum luctusquam ad domum convivii;in illa enim finis cunctorum hominum,et vivens hoc conferet in corde.
ECCL|7|3|Melior est tristitia risu,quia per tristitiam vultus corrigitur animus.
ECCL|7|4|Cor sapientium in domo luctus,et cor stultorum in domo laetitiae.
ECCL|7|5|Melius est a sapiente corripiquam laetari stultorum canticis,
ECCL|7|6|quia sicut sonitus spinarum ardentium sub olla,sic risus stulti.Sed et hoc vanitas.
ECCL|7|7|Quia calumnia stultum facit sapientem,et munus cor insanire facit.
ECCL|7|8|" Melior est finis negotii quam principium,melior est patiens arrogante ".
ECCL|7|9|Ne sis velox in animo ad irascendum, quia ira in sinu stulti requiescit.
ECCL|7|10|Ne dicas: "Quid, putas, causae est quod priora tempora meliora fuere quam nunc sunt? ". Non enim ex sapientia interrogas de hoc.
ECCL|7|11|Bona est sapientia cum divitiis et prodest videntibus solem.
ECCL|7|12|Sicut enim protegit sapientia, sic protegit pecunia; hoc autem plus habet eruditio, quod sapientia vitam tribuit possessori suo.
ECCL|7|13|Considera opera Dei: quod nemo possit corrigere, quod ille curvum fecerit.
ECCL|7|14|In die bona fruere bonis et in die mala considera: sicut hanc, sic et illam fecit Deus, ita ut non inveniat homo quidquam de futuro.
ECCL|7|15|Cuncta vidi in diebus vanitatis meae: est iustus, qui perit in iustitia sua, et impius, qui multo vivit tempore in malitia sua.
ECCL|7|16|Noli esse nimis iustusneque sapiens supra modum!Cur te perdere vis?
ECCL|7|17|Ne agas nimis impieet noli esse stultus!Cur mori debeas in tempore non tuo?
ECCL|7|18|Bonum est ut, quod habes, teneas, sed et ab illo ne subtrahas manum tuam, quia qui timet Deum, utrumque devitat.
ECCL|7|19|Sapientia confortabit sapientem super decem principes civitatis.
ECCL|7|20|Nullus enim homo iustus in terra, qui faciat bonum et non peccet.
ECCL|7|21|Sed et cunctis sermonibus, qui dicuntur, ne accommodes cor tuum, ne forte audias servum tuum maledicentem tibi;
ECCL|7|22|scit enim conscientia tua, quia et tu crebro maledixisti aliis.
ECCL|7|23|Cuncta tentavi in sapientia, dixi: " Sapiens efficiar ".
ECCL|7|24|Et ipsa longius recessit a me. Longe est, quod fuit; et alta est profunditas. Quis inveniet eam?
ECCL|7|25|Lustravi universa animo meo, ut scirem et considerarem et quaererem sapientiam et rationem et ut cognoscerem impietatem esse stultitiam et errorem imprudentiam.
ECCL|7|26|Et invenio amariorem morte mulierem, quae laqueus venatorum est, et sagena cor eius, vincula sunt manus illius. Qui placet Deo, effugiet eam; qui autem peccator est, capietur ab illa.
ECCL|7|27|Ecce hoc inveni, dixit Ecclesiastes, unum et alterum, ut invenirem rationem,
ECCL|7|28|quam adhuc quaerit anima mea, et non inveni:Hominem de mille unum repperi,mulierem ex omnibus non inveni.
ECCL|7|29|Ecce solummodo hoc inveni:Quod fecerit Deus hominem rectum,et ipsi quaesierint infinitas quaestiones.
ECCL|8|1|Quis talis, ut sapiens est?Et quis cognovit solutionem re rum?Sapientia hominis illuminat vultum eius,et durities faciei illius commutatur.
ECCL|8|2|Os regis observa et propter iuramenta Dei
ECCL|8|3|ne festines recedere a facie eius neque permaneas in re mala, quia omne, quod voluerit, faciet.
ECCL|8|4|Quia sermo illius potestate plenus est, nec dicere ei quisquam potest: " Quare ita facis? ".
ECCL|8|5|Qui custodit praeceptum, non experietur quidquam mali; tempus et iudicium cor sapientis intellegit.
ECCL|8|6|Omni enim negotio tempus est et iudicium, et multa hominis afflictio;
ECCL|8|7|ignorat enim quid futurum sit, nam quomodo sit futurum, quis nuntiabit ei?
ECCL|8|8|Non est in hominis potestate dominari super spiritum nec cohibere spiritum, nec habet potestatem supra diem mortis, nec ulla remissio est ingruente bello, neque salvabit impietas impium.
ECCL|8|9|Omnia haec consideravi et dedi cor meum cunctis operibus, quae fiunt sub sole, quo tempore dominatur homo homini in malum suum.
ECCL|8|10|Et ita vidi impios sepultos, discedentes de loco sancto; in oblivionem cadere in civitate, quod ita egerunt: sed et hoc vanitas est.
ECCL|8|11|Etenim, quia non profertur cito sententia contra opera mala, ideo cor filiorum hominum repletur, ut perpetrent mala.
ECCL|8|12|Nam peccator centies facit malum et prolongat sibi dies; verumtamen novi quod erit bonum timentibus Deum, qui verentur faciem eius.
ECCL|8|13|Non sit bonum impio, nec prolongabit dies suos quasi umbram, qui non timet faciem Domini.
ECCL|8|14|Est vanitas, quae fit super terram: sunt iusti, quibus mala proveniunt, quasi opera egerint impiorum, et sunt impii, quibus bona proveniunt, quasi iustorum facta habeant; sed et hoc vanissimum iudico.
ECCL|8|15|Laudavi igitur laetitiam quod non esset homini bonum sub sole, nisi quod comederet et biberet atque gauderet et hoc solum secum auferret de labore suo in diebus vitae suae, quos dedit ei Deus sub sole.
ECCL|8|16|Cum apposui cor meum, ut scirem sapientiam et intellegerem occupationem, quae versatur in terra, quod diebus et noctibus somnum non capit oculis,
ECCL|8|17|ecce intellexi quod omnium operum Dei nullam possit homo invenire rationem eorum, quae fiunt sub sole; et quanto plus laboraverit homo ad quaerendum, tanto minus inveniet; etiamsi dixerit sapiens se nosse, non poterit reperire.
ECCL|9|1|Omnia haec contuli in corde meo, ut curiose intellegerem quod iusti atque sapientes et opera eorum sunt in manu Dei. Utrum amor sit an odium, omnino nescit homo: coram illis omnia.
ECCL|9|2|Sicut omnibus sors una:iusto et impio,bono et malo,mundo et immundo,immolanti victimas et non immolanti.Sicut bonus sic et peccator;ut qui iurat, ita et ille qui iuramentum timet.
ECCL|9|3|Hoc est pessimum inter omnia, quae sub sole fiunt, quia sors eadem cunctis; unde et corda filiorum hominum implentur malitia et stultitia in vita sua, et novissima eorum apud mortuos.
ECCL|9|4|Qui enim sociatur omnibus viventibus, habet fiduciam: melior est canis vivus leone mortuo.
ECCL|9|5|Viventes enim sciunt se esse morituros; mortui vero nihil noverunt amplius nec habent ultra mercedem, quia oblivioni tradita est memoria eorum.
ECCL|9|6|Amor quoque eorum et odium et invidiae simul perierunt, nec iam habent partem in hoc saeculo et in opere, quod sub sole geritur.
ECCL|9|7|Vade ergo et comede in laetitia panem tuumet bibe cum gaudio vinum tuum,etenim iam diu placuerunt Deo opera tua.
ECCL|9|8|Omni tempore sint vestimenta tua candida,et oleum de capite tuo non deficiat.
ECCL|9|9|Perfruere vita cum uxore, quam diligis, cunctis diebus vitae instabilitatis tuae, qui dati sunt tibi sub sole omni tempore vanitatis tuae: haec est enim pars in vita et in labore tuo, quo laboras sub sole.
ECCL|9|10|Quodcumque facere potest manus tua, instanter operare, quia nec opus nec ratio nec sapientia nec scientia erunt apud inferos, quo tu properas.
ECCL|9|11|Verti me ad aliud et vidi sub sole nec velocium esse cursum nec fortium bellum nec sapientium panem nec doctorum divitias nec prudentium gratiam, sed tempus casumque in omnibus.
ECCL|9|12|Insuper nescit homo finem suum, sed sicut pisces capiuntur sagena mala, et sicut aves laqueo comprehenduntur, sic capiuntur homines in tempore malo, cum eis extemplo supervenerit.
ECCL|9|13|Hanc quoque sub sole vidi sapientiam et probavi maximam:
ECCL|9|14|civitas parva, et pauci in ea viri; venit contra eam rex magnus et vallavit eam exstruxitque munitiones magnas per gyrum.
ECCL|9|15|Inventusque est in ea vir pauper et sapiens et liberavit urbem per sapientiam suam; et nullus deinceps recordatus est hominis illius pauperis.
ECCL|9|16|Et dicebam ego meliorem esse sapientiam fortitudine,sed sapientia pauperis contemnitur,et verba eius non sunt audita.
ECCL|9|17|Verba sapientium cum lenitate audiunturplus quam clamor principis inter stultos.
ECCL|9|18|Melior est sapientia quam arma bellica;sed unus, qui peccaverit, multa bona perdet.
ECCL|10|1|Muscae morientes perdunt et corrumpunt oleum unguentarii.Gravior quam sapientia et gloria est parva stultitia.
ECCL|10|2|Cor sapientis in dextera eius,et cor stulti in sinistra illius.
ECCL|10|3|Sed et in via stultus ambulans, cum ipse insipiens sit, omnes stultos aestimat.
ECCL|10|4|Si spiritus potestatem habentis ascenderit contra te, locum tuum ne dimiseris, quia lenitas faciet cessare peccata maxima.
ECCL|10|5|Est malum, quod vidi sub sole quasi errorem egredientem a facie principis:
ECCL|10|6|positum stultum in dignitate sublimi et divites sedere deorsum.
ECCL|10|7|Vidi servos in equis et principes ambulantes super terram quasi servos.
ECCL|10|8|Qui fodit foveam, incidet in eam;et, qui dissipat murum, mordebit eum coluber.
ECCL|10|9|Qui excidit lapides, affligetur in eis;et, qui scindit ligna, periclitabitur ex eis.
ECCL|10|10|Si retusum fuerit ferrum, et aciem eius non exacueris, labor multiplicabitur, sed lucrum industriae erit sapientia.
ECCL|10|11|Si mordeat serpens incantatione neglecta, nihil lucri habet incantator.
ECCL|10|12|Verba oris sapientis gratia,et labia insipientis praecipitabunt eum.
ECCL|10|13|Initium verborum eius stultitia,et novissimum oris illius insipientia mala.
ECCL|10|14|Stultus verba multiplicat: Ignorat homo quid futurum sit;et, quid post se futurum sit, quis ei poterit indicare?".
ECCL|10|15|Labor stultorum affliget eos,qui nesciunt in urbem pergere.
ECCL|10|16|Vae tibi, terra, cuius rex puer est,et cuius principes mane comedunt.
ECCL|10|17|Beata terra, cuius rex nobilis est,et cuius principes vescuntur in tempore suoad reficiendum et non ad luxuriam.
ECCL|10|18|In pigris manibus humiliabitur contignatio,et in remissis perstillabit domus.
ECCL|10|19|In risum faciunt epulas;vinum laetificat vitam,et pecunia praestat omnia.
ECCL|10|20|In cogitatione tua regi ne detrahaset in secreto cubiculi tui ne maledixeris diviti,quia et aves caeli portabunt vocem tuam,et, qui habet pennas, annuntiabit sententiam.
ECCL|11|1|Mitte panem tuum super transeuntes aquas, quia post tempora multa invenies illum.
ECCL|11|2|Da partem septem necnon et octo, quia ignoras, quid futurum sit mali super terram.
ECCL|11|3|Si repletae fuerint nubes,imbrem super terram effundent;si ceciderit lignum ad austrum aut ad aquilonem,in quocumque loco ceciderit, ibi erit.
ECCL|11|4|Qui observat ventum, non seminat, et, qui considerat nubes, numquam metet.
ECCL|11|5|Quomodo ignoras, quae sit via spiritus, et qua ratione compingantur ossa in ventre praegnantis, sic nescis opera Dei, qui fabricator est omnium.
ECCL|11|6|Mane semina semen tuum,et vespere ne cesset manus tua,quia nescis quid magis prosit,hoc aut illud,et si utrumque simul melius erit.
ECCL|11|7|Dulce lumen,et delectabile est oculis videre solem.
ECCL|11|8|Si annis multis vixerit homoet in his omnibus laetatus fuerit,meminisse debet tenebrosi temporis, quod multum erit:omne, quod venerit, vanitas.
ECCL|11|9|Laetare ergo, iuvenis, in adulescentia tua,et in bono sit cor tuum in diebus iuventutis tuae,et ambula in viis cordis tuiet in intuitu oculorum tuorumet scito quod pro omnibus hisadducet te Deus in iudicium.
ECCL|11|10|Aufer curam a corde tuoet amove malum a carne tua;adulescentia enim et iuventus vanae sunt.
ECCL|12|1|Memento Creatoris tuiin diebus iuventutis tuae,antequam veniat tempus afflictionis,et appropinquent anni, de quibus dicas: Non mihi placent ";
ECCL|12|2|antequam tenebrescatsol et lumen et luna et stellae,et revertantur nubes post pluviam;
ECCL|12|3|quando commovebuntur custodes domus,et nutabunt viri fortissimi,et otiosae erunt molentes imminuto numero,et tenebrescent videntes per foramina,
ECCL|12|4|et claudentur ostia in plateasubmissa voce molentis,et consurgent ad vocem volucris,et subsident omnes filiae carminis;
ECCL|12|5|excelsa quoque timebuntet formidabunt in via.Florebit amygdalus,reptabit locusta,et dissipabitur capparis,quoniam ibit homo in domum aeternitatis suae,et circuibunt in platea plangentes,
ECCL|12|6|antequam rumpatur funiculus argenteus,et frangatur lecythus aureus,et conteratur hydria super fontem,et confringatur rota super cisternam,
ECCL|12|7|et revertatur pulvis in terram suam, unde erat,et spiritus redeat ad Deum, qui dedit illum.
ECCL|12|8|Vanitas vanitatum,dixit Ecclesiastes,et omnia vanitas.
ECCL|12|9|Cumque esset sapientissimus, Ecclesiastes docuit insuper populum scientiam; ponderavit et investigans composuit parabolas multas.
ECCL|12|10|Quaesivit Ecclesiastes verba delectabilia et conscripsit sermones rectissimos ac veritate plenos.
ECCL|12|11|Verba sapientium sicut stimuli, et quasi clavi defixi sunt magistri collationum; data sunt a pastore uno.
ECCL|12|12|His amplius, fili mi, ne requiras: faciendi plures libros nullus est finis, frequensque meditatio carnis afflictio est.
ECCL|12|13|Finis loquendi, omnibus auditis: Deum time et mandata eius observa; hoc est enim omnis homo.
ECCL|12|14|Et cuncta, quae fiunt, adducet Deus in iudicium circa omne occultum, sive bonum sive malum.
