ZECH|1|1|大流士 王第二年八月，耶和华的话临到 易多 的孙子， 比利家 的儿子 撒迦利亚 先知，说：
ZECH|1|2|“耶和华曾向你们祖先大发烈怒。
ZECH|1|3|你要对 以色列 人说，万军之耶和华如此说：你们要转向我，这是万军之耶和华说的，我就转向你们，这是万军之耶和华说的。
ZECH|1|4|不要效法你们的祖先。从前的先知呼叫他们说：‘万军之耶和华如此说，当回转离开你们的恶道恶行。’他们却不听，也不顺从我。这是耶和华说的。
ZECH|1|5|你们的祖先在哪里呢？那些先知能永远存活吗？
ZECH|1|6|然而我的言语和律例，就是我所吩咐我仆人众先知的，岂不临到你们的祖先吗？他们就回转，说：万军之耶和华定意按我们的所作所为对待我们，他也已经照样行了。”
ZECH|1|7|大流士 第二年十一月，就是细罢特月二十四日，耶和华的话临到 易多 的孙子， 比利家 的儿子 撒迦利亚 先知，说：
ZECH|1|8|“我夜间观看，看哪，有一人骑着红马，站在洼地的番石榴树中间。在他身后有红色、褐色和白色的马。”
ZECH|1|9|我说：“主啊，这是什么意思？”与我说话的天使说：“我要指示你这是什么意思。”
ZECH|1|10|那站在番石榴树中间的人回答说：“这是奉耶和华差遣，在遍地巡逻的。”
ZECH|1|11|他们对站在番石榴树中间耶和华的使者说：“我们在遍地巡逻，看哪，全地都安息平静。”
ZECH|1|12|于是，耶和华的使者说：“万军之耶和华啊，你恼恨 耶路撒冷 和 犹大 的城镇已经七十年了，你不施怜悯要到几时呢？”
ZECH|1|13|耶和华就用美善的话和安慰的话回答那与我说话的天使。
ZECH|1|14|与我说话的天使对我说：“你要宣告，万军之耶和华如此说：我为 耶路撒冷 而妒忌，为 锡安 大大妒忌。
ZECH|1|15|我非常恼怒那享安逸的列国，因我从前稍微恼怒，他们就越发加害。
ZECH|1|16|所以耶和华如此说：现在我回到 耶路撒冷 ，仍要施怜悯，我的殿要重建在其中，准绳必拉在 耶路撒冷 之上。这是万军之耶和华说的。
ZECH|1|17|你要再宣告，万军之耶和华如此说：我的城镇要再度繁荣发达。耶和华必再安慰 锡安 ，拣选 耶路撒冷 。”
ZECH|1|18|我举目观看，看哪，有四只角。
ZECH|1|19|我问那与我说话的天使：“这是什么意思？”他对我说：“这是击散 犹大 、 以色列 和 耶路撒冷 的角。”
ZECH|1|20|耶和华又把四个匠人指给我看。
ZECH|1|21|我问：“这些人来做什么呢？”他说：“那是击散 犹大 的角，使人不敢抬头；但这些匠人前来威吓列国，打掉列国的角，因为他们举起角来击散 犹大 地。”
ZECH|2|1|我举目观看，看哪，有一人手拿丈量的绳。
ZECH|2|2|我问：“你到哪里去？”他对我说：“要去丈量 耶路撒冷 ，看有多宽多长。”
ZECH|2|3|看哪，与我说话的天使出去 ，另有一位天使迎着他来，
ZECH|2|4|对他说：“你跑去告诉这个年轻人说， 耶路撒冷 必有人居住，如同无城墙的乡村，因为其中的人和牲畜很多。
ZECH|2|5|耶和华说：‘我要作 耶路撒冷 四围火的城墙，并要作城中的荣耀。’”
ZECH|2|6|耶和华说：“来，来！你们要从北方之地逃回；因我曾把你们分散到天的四方 。这是耶和华说的。”
ZECH|2|7|来！住 巴比伦 的 锡安 百姓啊，逃吧！
ZECH|2|8|万军之耶和华在显出荣耀之后，差遣我到掳掠你们的列国那里，他如此说：“碰你们的就是碰他自己 眼中的瞳人。
ZECH|2|9|看哪，我要挥手攻击他们，他们就必作自己奴仆的掳物。”你们就知道万军之耶和华差遣了我。
ZECH|2|10|耶和华说：“ 锡安 哪，应当欢乐歌唱，因为，看哪，我要来，要住在你中间。
ZECH|2|11|在那日，必有许多国家归附耶和华，作我的子民。我要住 在你中间。”你就知道万军之耶和华差遣我到你那里去。
ZECH|2|12|耶和华必收回 犹大 ，作为他圣地的产业，他必再度拣选 耶路撒冷 。
ZECH|2|13|凡血肉之躯都当在耶和华面前静默无声，因为他从他的圣所奋起了。
ZECH|3|1|天使 指给我看： 约书亚 大祭司站在耶和华的使者面前，撒但站在 约书亚 的右边控告他。
ZECH|3|2|耶和华向撒但说：“撒但哪，耶和华责备你！拣选 耶路撒冷 的耶和华责备你！这不是从火中抽出来的一根柴吗？”
ZECH|3|3|约书亚 穿着污秽的衣服，站在那使者面前。
ZECH|3|4|使者吩咐那些侍立在他面前的说：“脱去他污秽的衣服。”又对 约书亚 说：“你看，我使你的罪孽离开你，要给你穿上华美的衣服。”
ZECH|3|5|我说 ：“要将洁净的冠冕戴在他头上。”他们就把洁净的冠冕戴在他头上，给他穿上华美的衣服，耶和华的使者在旁边站立。
ZECH|3|6|耶和华的使者告诫 约书亚 说，
ZECH|3|7|万军之耶和华如此说：“你若遵行我的道，谨守我的命令，就可以管理我的家，看守我的院宇；我也要使你在这些侍立的人中间来往。
ZECH|3|8|约书亚 大祭司啊，你和坐在你面前的同伴都当听，因为他们是作预兆的：看哪，我必使我仆人 大卫 的苗裔 长出。
ZECH|3|9|看哪，这是我在 约书亚 面前所立的石头，这一块石头上有七眼。看哪，我要亲自雕刻这石头，并在一日之间除掉这地的罪孽。这是万军之耶和华说的。
ZECH|3|10|在那日，你们各人要请邻舍坐在葡萄树和无花果树下。这是万军之耶和华说的。”
ZECH|4|1|那与我说话的天使又来叫醒我，好像人睡觉时被唤醒一样。
ZECH|4|2|他问我：“你看见什么？”我说：“我看见了，看哪，有一个纯金的灯台，顶上有灯座，其上有七盏灯，每盏灯的上头有七根管子；
ZECH|4|3|旁边有两棵橄榄树，一棵在灯座的右边，一棵在灯座的左边。”
ZECH|4|4|我问与我说话的天使说：“主啊，这是什么意思？”
ZECH|4|5|与我说话的天使回答，对我说：“你不知道这是什么意思吗？”我说：“主啊，我不知道。”
ZECH|4|6|他回答我说：“这是耶和华指示 所罗巴伯 的话。万军之耶和华说：不是倚靠势力，不是倚靠才能，乃是倚靠我的灵方能成事 。
ZECH|4|7|大山哪，你算什么呢？在 所罗巴伯 面前，你必夷为平地。他安放顶上的那块石头，人就欢呼：‘愿恩惠、恩惠归与这殿！’”
ZECH|4|8|耶和华的话临到我，说：
ZECH|4|9|“ 所罗巴伯 的手立了这殿的根基，他的手也必完成这工，你就知道万军之耶和华差遣我到你们这里。
ZECH|4|10|谁藐视这日的事为小呢？他们见 所罗巴伯 手拿石垂线就欢喜。这七盏灯 是耶和华的眼睛，遍察全地。”
ZECH|4|11|我问天使说：“那么在灯台左右的这两棵橄榄树是什么意思呢？”
ZECH|4|12|我再次问他：“这两根橄榄树枝在两根流出金色油的金嘴旁边，是什么意思呢？”
ZECH|4|13|他对我说：“你不知道这是什么意思吗？”我说：“主啊，我不知道。”
ZECH|4|14|他说：“这是两位受膏者，侍立在全地之主的旁边。”
ZECH|5|1|我又举目观看，看哪，有一飞行的书卷。
ZECH|5|2|他问我：“你看见什么？”我回答：“我看见一飞行的书卷，长二十肘，宽十肘。”
ZECH|5|3|他对我说：“这就是向全地面发出的诅咒。凡偷窃的必按书卷这面的话除灭，凡起假誓的必按书卷那面的话除灭。
ZECH|5|4|万军之耶和华说：我要把这书卷送出去，进入偷窃者的家和指着我名起假誓者的家，停留在他家里，连房屋带木头和石头都毁灭了。”
ZECH|5|5|与我说话的天使前来，对我说：“你要举目观看，看那出现的是什么。”
ZECH|5|6|我问：“这是什么呢？”他说：“这出现的是量器 。”又说：“是他们的眼目，遍行全地 。”
ZECH|5|7|看哪，圆形的铅盖被抬起来，有一个妇人坐在量器中。
ZECH|5|8|天使说：“这是罪恶。”他就把妇人推进量器里，把铅盖压在量器的口上。
ZECH|5|9|于是我举目观看，看哪，有两个妇人前来，她们的翅膀中有风，翅膀如同鹳鸟的翅膀。她们把量器抬起来，悬在天地之间。
ZECH|5|10|我问那与我说话的天使：“她们要把量器抬到哪里去呢？”
ZECH|5|11|他对我说：“要抬到 示拿 地去，为它建造房屋；等预备妥当，就把它安放在自己的台座上。”
ZECH|6|1|我又举目观看，看哪，有四辆马车从两座山的中间出来；那两座山是铜山。
ZECH|6|2|第一辆车套着红马，第二辆车套着黑马，
ZECH|6|3|第三辆车套着白马，第四辆车套着带斑点的马，都是强壮的 。
ZECH|6|4|我就回应与我说话的天使说：“主啊，这是什么意思？”
ZECH|6|5|天使回答，对我说：“这是天的四风，是从全地之主面前出来的。”
ZECH|6|6|套着黑马的车往北方之地去，白马跟随在后；有斑点的马往南方之地去；
ZECH|6|7|那些壮马出来，急着要在地上巡逻。天使说：“你们只管在地上巡逻。”它们就在地上巡逻。
ZECH|6|8|他又呼叫我，告诉我说：“你看，往北方地去的已在北方之地使我放心。”
ZECH|6|9|耶和华的话临到我，说：
ZECH|6|10|“你要拿从 巴比伦 归来的被掳之人 黑玳 、 多比雅 、 耶大雅 所献的，当日就要进到 西番雅 的儿子 约西亚 的家里，
ZECH|6|11|拿这金银做冠冕，戴在 约撒答 的儿子 约书亚 大祭司的头上；
ZECH|6|12|对他说，万军之耶和华如此说：‘看哪，那名称为 大卫 苗裔的，要在本处生长，并要建造耶和华的殿。
ZECH|6|13|就是他，要建造耶和华的殿，他要承受尊荣，坐在位上掌王权；又有一位祭司坐在自己的位上，两职之间筹划和平。
ZECH|6|14|这冠冕要归 希连 、 多比雅 、 耶大雅 ，和 西番雅 的儿子 贤 ，放在耶和华的殿里作为纪念。’”
ZECH|6|15|远方的人要来建造耶和华的殿，你们因此就知道，万军之耶和华差遣我到你们这里来。你们若留意听从耶和华－你们上帝的话，这事必然成就。
ZECH|7|1|大流士 王第四年九月，就是基斯流月初四，耶和华的话临到 撒迦利亚 。
ZECH|7|2|那时 伯特利 人已经差遣 沙利色 和 利坚．米勒 ，并他们的人，去恳求耶和华的恩，
ZECH|7|3|问万军之耶和华殿中的祭司，又问先知：“我当如历年以来所行，在五月哭泣斋戒吗？”
ZECH|7|4|万军之耶和华的话临到我，说：
ZECH|7|5|“你要向这地全体百姓和祭司说：‘你们这七十年来，在五月、七月禁食悲哀，岂是真的向我禁食吗？
ZECH|7|6|你们吃喝，不是为自己吃，为自己喝吗？
ZECH|7|7|当 耶路撒冷 和四围的城镇有人居住，享繁荣， 尼革夫 和 谢非拉 也有人居住的时候，耶和华藉从前的先知所宣告的，你们不当听吗？’”
ZECH|7|8|耶和华的话临到 撒迦利亚 ，说：
ZECH|7|9|“万军之耶和华如此说：你们要按真正的公平来审判，彼此以慈爱怜悯相待。
ZECH|7|10|不可欺压寡妇、孤儿、寄居的和困苦的人。谁都不可心里谋害弟兄。
ZECH|7|11|他们却不留意；耸肩悖逆，耳朵发沉，不肯听从。
ZECH|7|12|他们的心坚硬如金刚石，不听律法和万军之耶和华藉着他的灵差遣从前先知所说的话。因此，万军之耶和华大发烈怒。
ZECH|7|13|万军之耶和华说：我曾呼唤他们，他们不听；将来他们呼求我，我也不听！
ZECH|7|14|我必以旋风将他们吹散到素不认识的万国中。他们离开以后，地就荒凉，无人来往经过；他们使美好之地荒凉了。”
ZECH|8|1|万军之耶和华的话临到我，说：
ZECH|8|2|“万军之耶和华如此说：我为 锡安 而妒忌，大大妒忌；我为了它妒忌而大发烈怒。
ZECH|8|3|耶和华如此说：我要回到 锡安 ，住在 耶路撒冷 中间。 耶路撒冷 必称为忠实的城，万军之耶和华的山必称为圣山。
ZECH|8|4|万军之耶和华如此说：将来必有年老的男女坐在 耶路撒冷 的广场上，各人因年纪老迈而手拿枴杖。
ZECH|8|5|城里的广场满有男孩女孩在玩耍。
ZECH|8|6|万军之耶和华如此说：在那些日子，即使这事在这余民眼中看为奇妙，难道在我眼中也看为奇妙吗？这是万军之耶和华说的。
ZECH|8|7|万军之耶和华如此说：看哪，我要从日出之地、从日落之地拯救我的子民。
ZECH|8|8|我要领他们来，使他们住在 耶路撒冷 中间。他们要作我的子民，我要作他们的上帝，都凭信实和公义。
ZECH|8|9|“万军之耶和华如此说：你们的手要坚强；这些日子，你们已听见先知的口，在万军之耶和华殿的根基立定、圣殿建造的日子所说的这些话。
ZECH|8|10|那些日子以前，人得不着工价，牲畜也无人雇用；且因敌人的缘故，出入不得平安；因我使人与人互相攻击。
ZECH|8|11|但如今，我对这余民必不像先前的日子。这是万军之耶和华说的。
ZECH|8|12|因为他们要平安撒种，葡萄树要结果子，土地必有出产，天也必降甘露。我要使这余民享受这一切。
ZECH|8|13|犹大 家和 以色列 家啊，你们从前在列国中怎样成为可诅咒的；照样，我要拯救你们，使你们得福 。不要惧怕，你们的手要坚强。
ZECH|8|14|“万军之耶和华如此说：你们祖先惹我发怒的时候，我怎样定意降祸，并不改变；万军之耶和华说，
ZECH|8|15|这些日子我也定意施恩给 耶路撒冷 和 犹大 家；你们不要惧怕。
ZECH|8|16|你们所当行的是这样：每个人要与邻舍说诚实话，在城门口要按真正的公平来审判，使人和睦。
ZECH|8|17|谁都不可心里谋害邻舍，也不可喜爱起假誓，因为这些事都为我所恨恶。这是耶和华说的。”
ZECH|8|18|万军之耶和华的话临到我，说：
ZECH|8|19|“万军之耶和华如此说：四月的禁食、五月的禁食、七月的禁食和十月的禁食，必成为 犹大 家的欢喜和快乐，以及美好的节期；所以你们要喜爱诚实与和平。
ZECH|8|20|“万军之耶和华如此说：将来还有众百姓和许多城镇的居民要来。
ZECH|8|21|这城的居民必到那城，说：‘我们快去恳求耶和华的恩，寻求万军之耶和华；我自己也要去。’
ZECH|8|22|必有许多民族和强盛的国家来到 耶路撒冷 寻求万军之耶和华，恳求耶和华的恩。
ZECH|8|23|万军之耶和华如此说：在那些日子，列国中说各种语言的人，必有十个人强拉住一个 犹大 人衣服的边，说：‘我们要与你们同去，因为我们听见上帝与你们同在了。’”
ZECH|9|1|耶和华的默示， 他的话临到 哈得拉 地、 大马士革 －因世人和 以色列 各支派的眼目都向着耶和华－
ZECH|9|2|和邻近的 哈马 ， 以及 推罗 和 西顿 。 因为它极有智慧，
ZECH|9|3|推罗 为自己建造坚固城 ， 堆起银子如尘沙， 纯金如街上的泥土。
ZECH|9|4|看哪，主必赶出它， 重创它海上的势力， 它必被火吞灭。
ZECH|9|5|亚实基伦 看见必惧怕， 迦萨 看见甚痛苦， 以革伦 因失了盼望而蒙羞； 迦萨 必不再有君王， 亚实基伦 也不再有人居住，
ZECH|9|6|混血的人要住在 亚实突 ； 我必除灭 非利士 人的骄傲。
ZECH|9|7|我要除去他口中带血之肉 和牙齿内可憎之物。 他必作余民归于我们的上帝， 在 犹大 像族长一样； 以革伦 必如 耶布斯 人。
ZECH|9|8|我要扎营在我的家， 敌军不得任意往来， 暴虐的人也不再经过， 因为我亲眼看顾。
ZECH|9|9|锡安 哪，应当大大喜乐； 耶路撒冷 啊，应当欢呼。 看哪，你的王来到你这里！ 他是公义的，并且施行拯救， 谦和地骑着驴， 骑着小驴，驴的驹子。
ZECH|9|10|我必除灭 以法莲 的战车 和 耶路撒冷 的战马； 战争的弓也必剪除。 他要向列国讲和平； 他的权柄必从这海管到那海， 从 大河 管到地极。
ZECH|9|11|锡安 哪，我因与你立约的血， 要从无水坑里释放你中间被囚的人。
ZECH|9|12|被囚而有指望的人哪，要转回堡垒； 我今日宣告，我必加倍补偿你。
ZECH|9|13|我为自己把 犹大 弯紧， 我使 以法莲 如满弓。 锡安 哪，我要唤起你的儿女， 希腊 啊，我要攻击你的儿女， 使你如勇士的刀。
ZECH|9|14|耶和华要显现在他们身上， 他的箭要射出如闪电。 主耶和华必吹角， 乘南方的旋风而行。
ZECH|9|15|万军之耶和华必保护他们； 他们要吞灭，要践踏弹弓的石头 ； 他们呐喊，狂饮 如喝酒， 如盛满的碗， 又如坛的四角。
ZECH|9|16|当那日，耶和华－他们的上帝 必看他的百姓如羊群，拯救他们； 因为他们如冠冕上的宝石， 在他的地上如旗帜高举 。
ZECH|9|17|他是何等善！ 他是何其美！ 五谷使少男强壮， 新酒使少女健美。
ZECH|10|1|春雨的季节，你们要向耶和华求雨。 耶和华发出雷电， 为众人降下大雨， 把田园的菜蔬赐给人。
ZECH|10|2|因为家中神像所言的是虚空， 占卜者所见的是虚假， 他们讲说假梦， 徒然安慰人。 所以众人如羊流离， 因无牧人就受欺压。
ZECH|10|3|我的怒气向牧人发作， 我必惩罚那为首的 ； 万军之耶和华眷顾他的羊群， 就是 犹大 家， 必使他们如战场上的骏马。
ZECH|10|4|房角石从他而出， 橛子从他而出， 战争的弓也从他而出， 每一个掌权的都从他而出。
ZECH|10|5|他们必如战场上的勇士， 践踏仇敌如街上的泥土。 他们必争战，因为耶和华与他们同在， 他们必使骑马的羞愧。
ZECH|10|6|我要坚固 犹大 家， 拯救 约瑟 家， 我要领他们归回，因我怜悯他们， 他们必像我未曾弃绝他们一样； 都因我是耶和华－他们的上帝， 我必应允他们。
ZECH|10|7|以法莲 人必如勇士， 他们心中畅快如同喝酒； 他们的儿女看见就欢喜， 他们的心必因耶和华喜乐。
ZECH|10|8|我要呼叫，聚集他们， 因我已经救赎他们。 他们的人数必增添， 如从前增添一样。
ZECH|10|9|我要将他们分散在列国中， 他们必在远方记得我； 他们与儿女都必存活， 他们要归回。
ZECH|10|10|我必使他们从 埃及 地归回， 从 亚述 召集他们， 领他们到 基列 地和 黎巴嫩 ； 这些还不够他们居住。
ZECH|10|11|耶和华 必经过苦海，击打海浪。 尼罗河 的深处全都枯干， 亚述 的骄傲必降卑， 埃及 的权杖必除去。
ZECH|10|12|我要使他们倚靠耶和华，得以坚固， 他们必奉他的名而行 ； 这是耶和华说的。
ZECH|11|1|黎巴嫩 哪，敞开你的门， 任火吞灭你的香柏树。
ZECH|11|2|哀号吧，松树！ 因为香柏树倾倒了，高大的树毁坏了。 哀号吧， 巴珊 的橡树！ 因为茂盛的树林倒下来了。
ZECH|11|3|听啊，有牧人在哀号， 因他们的荣华败落了； 听啊，有少壮狮子咆哮， 因 约旦河 旁的丛林荒废了。
ZECH|11|4|耶和华－我的上帝如此说：“你要牧养这群将宰的羊。
ZECH|11|5|买羊的宰了他们，却不认为自己有罪；卖他们的也说：‘耶和华是应当称颂的，因我富足了。’牧养他们的并不怜悯他们。
ZECH|11|6|我不再怜悯这地的居民。看哪，我要将这些人交在各人的邻舍和君王手中；他们必毁灭这地，我却不救任何一个脱离他们的手。这是耶和华说的。”
ZECH|11|7|于是，我牧养这群将宰的羊，就是羊群中最困苦的 ；我拿着两根杖，一根我称为“恩惠” ，一根称为“联合”。这样，我就牧养这群羊。
ZECH|11|8|一个月之内，我废除了三个牧人，因为我的心厌烦他们，他们的心也憎恶我。
ZECH|11|9|我就说：“我不牧养你们。要死的，由他死；灭亡的，由他灭亡；剩余的，由他们彼此吞食。”
ZECH|11|10|我拿起那根称为“恩惠”的杖，折断它，表明我废弃与万民所立的约。
ZECH|11|11|当日约就废了。因此，那些羊群中最困苦的 ，看着我，就知道这真是耶和华的话。
ZECH|11|12|我对他们说：“你们若看为美，就给我工价。不然，就罢了！”于是他们秤了三十块银钱作为我的工价。
ZECH|11|13|耶和华对我说：“把它丢给窑户。那是他们对我所估定的好价钱！”我就取这三十块银钱，在耶和华的殿中将它丢给窑户。
ZECH|11|14|我又折断第二根杖，就是称为“联合”的那根杖，表明我废弃 犹大 与 以色列 弟兄间的情谊。
ZECH|11|15|耶和华对我说：“你再把愚昧牧人所用的器具拿来，
ZECH|11|16|因为，看哪，我要在这地立一个牧人；他不看顾将亡的，不寻找分散的，不医治受伤的，也不牧养强壮的；却要吞吃肥羊的肉，撕裂它们的蹄。
ZECH|11|17|祸哉！无用的牧人丢弃羊群， 刀必临到他的膀臂和右眼上； 他的膀臂必全然枯干， 他的右眼也必昏暗失明。”
ZECH|12|1|耶和华的默示，他的话论到 以色列 。 铺张诸天、建立地基、造人里面之灵的耶和华说：
ZECH|12|2|“看哪，我要使 耶路撒冷 成为令四围列国百姓昏醉的杯； 耶路撒冷 被围困， 犹大 也一样受困 。
ZECH|12|3|在那日，我要使 耶路撒冷 成为万民的一块沉重石头，凡举起它的必受重伤；地上的万国都聚集攻击它。
ZECH|12|4|到那日，我必令一切的马匹惊惶，使骑马的癫狂。我必张开眼睛看顾 犹大 家，却使列国一切的马匹瞎眼。这是耶和华说的。
ZECH|12|5|犹大 的族长心里要说：‘ 耶路撒冷 的居民因倚靠万军之耶和华－他们的上帝，就成为我的力量 。’
ZECH|12|6|“那日，我必使 犹大 的族长如柴堆中的火盆，又如禾捆里的火把；他们必左右吞灭四围列国的百姓。 耶路撒冷 却仍屹立在本处，仍在 耶路撒冷 ！
ZECH|12|7|“耶和华要先拯救 犹大 的帐棚，免得 大卫 家的荣耀和 耶路撒冷 居民的荣耀胜过 犹大 。
ZECH|12|8|那日，耶和华必保护 耶路撒冷 的居民。他们中间软弱的在那日必如 大卫 ； 大卫 家必如上帝，如行在他们前面的耶和华的使者。
ZECH|12|9|那日，我必定意灭绝前来攻击 耶路撒冷 的万国。”
ZECH|12|10|“我要将那施恩与恳求的灵，浇灌 大卫 家和 耶路撒冷 的居民。他们必仰望我，就是他们所扎的那位。他们必为他悲伤，如丧独子，又为他哀哭，如丧长子。
ZECH|12|11|那日，在 耶路撒冷 必有大大的哀号，如 米吉多 平原上 哈达．临门 的哀号。
ZECH|12|12|这地必哀哭：一家一家地哭， 大卫 家的家族聚在一处，他们的妇女聚在一处； 拿单 家的家族聚在一处，他们的妇女聚在一处。
ZECH|12|13|利未 家的家族聚在一处，他们的妇女聚在一处； 示每 家的家族聚在一处，他们的妇女聚在一处。
ZECH|12|14|其余的各家，每一家的家族聚在一处，他们的妇女聚在一处。”
ZECH|13|1|“在那日，因罪恶与污秽的缘故，必有一泉源为 大卫 家和 耶路撒冷 的居民而开。”
ZECH|13|2|万军之耶和华说：“在那日，我要从地上除灭偶像的名，使它不再被记得；我也必使这地不再有先知，不再有污秽的灵。
ZECH|13|3|若还有人说预言，生他的父母必对他说：‘你不得存活，因为你假借耶和华的名说谎话。’生他的父母在他说预言时，要将他刺死。
ZECH|13|4|那日，凡作先知说预言的必因所论的异象羞愧，不再穿毛皮外袍哄骗人。
ZECH|13|5|他要说：‘我不是先知，我是耕地的；我从幼年就作人的奴仆。’
ZECH|13|6|有人对他说：‘你两手臂间是什么伤呢？’他说：‘这是我在亲友家中所受的伤。’”
ZECH|13|7|万军之耶和华说： 刀剑哪，兴起攻击我的牧人， 攻击我的同伴吧！ 要击打牧人，羊就分散了； 我必反手攻击那微小的。
ZECH|13|8|这全地的人， 三分之二将被剪除而死， 三分之一仍必存留。 这是耶和华说的。
ZECH|13|9|我要使这三分之一经过火， 熬炼他们，如熬炼银子； 试炼他们，如试炼金子。 他们要求告我的名， 我必应允他们。 我说：“这是我的子民。” 他们要说：“耶和华是我的上帝。”
ZECH|14|1|看哪，耶和华的日子临近了，你的财物必被抢掠，在你中间被瓜分。
ZECH|14|2|我要招聚万国与 耶路撒冷 争战；城必被攻取，房屋被抢夺，妇女被玷污，城中的一半被掳去；但其余的百姓不会从城中被剪除。
ZECH|14|3|那时，耶和华要出去与那些国家打仗，如同从前战争的日子打仗一样。
ZECH|14|4|那日，他的脚必站在 橄榄山 上，这山面向 耶路撒冷 的东边。 橄榄山 必从中间裂开，自东至西成为极大的谷；山的一半向北挪移，一半向南挪移。
ZECH|14|5|你们要从我的山谷中逃跑，因为山谷必延到 亚萨 。你们要逃跑，如在 犹大 王 乌西雅 年间逃避大地震一样 。耶和华－我的上帝必降临，所有的圣者与你 同来。
ZECH|14|6|在那日，必没有光，不会放晴，只有乌云 。
ZECH|14|7|耶和华所知道的那一日，没有白天，没有黑夜，到了晚上仍有亮光。
ZECH|14|8|在那日，必有活水从 耶路撒冷 出来，一半往东海流，一半往西海流；冬夏都是如此。
ZECH|14|9|耶和华要作全地的王。那日，耶和华必为独一无二，他的名也是独一无二。
ZECH|14|10|从 迦巴 直到 耶路撒冷 南方的 临门 ，全地要变为旷野。 耶路撒冷 要矗立于本处，从 便雅悯门 到 旧门 ，又到 角门 ，并从 哈楠业楼 ，直到王的酒池。
ZECH|14|11|人要住在其中，不再有诅咒； 耶路撒冷 必安然屹立。
ZECH|14|12|这是耶和华所降的灾殃，要攻击那些与 耶路撒冷 作战的万民；他们两脚站立时，肉要溃烂，眼在眶中溃烂，舌在口中也溃烂。
ZECH|14|13|那日，耶和华必使他们大大混乱。他们彼此用手揪住，用手互相攻击。
ZECH|14|14|犹大 也要在 耶路撒冷 打仗 。那时四围各国的财物，就是许许多多的金银和衣服，必被收聚。
ZECH|14|15|马匹、骡子、骆驼、驴和营中一切的牲畜所遭的灾殃与那灾殃一样。
ZECH|14|16|上来攻击 耶路撒冷 的列国中所有剩下的人，要年年上来敬拜大君王－万军之耶和华，并守住棚节。
ZECH|14|17|地上万族中，凡不上 耶路撒冷 敬拜大君王－万军之耶和华的，雨必不降在他们的地上。
ZECH|14|18|埃及 族若不上来，雨必不降在他们的地上；凡不上来守住棚节的列国，耶和华必用这灾攻击他们。
ZECH|14|19|这就是 埃及 的惩罚和那些不上来守住棚节之列国的惩罚。
ZECH|14|20|在那日，马的铃铛上要刻上“归耶和华为圣”。耶和华殿内的锅必如祭坛前的碗一样。
ZECH|14|21|耶路撒冷 和 犹大 一切的锅都必归万军之耶和华为圣。凡献祭的都必来取这锅，在其中煮肉。当那日，在万军之耶和华的殿中必不再有做买卖的人 。
