JER|1|1|Слова Єремії, сина Хілкійїного, з священиків, що в Анатоті, у Веніяминовому краї,
JER|1|2|що було до нього Господнє слово за днів Йосії, Амонового сина, Юдиного царя, тринадцятого року його царювання.
JER|1|3|І було воно й за днів Єгоякима, сина Йосіїного, Юдиного царя, аж до кінця одинадцятого року Седекії, сина Йосіїного, Юдиного царя, аж до виходу Єрусалиму на вигнання в п'ятому місяці.
JER|1|4|І прийшло мені слово Господнє, говорячи:
JER|1|5|Ще поки тебе вформував в утробі матерній, Я пізнав був тебе, і ще поки ти вийшов із нутра, тебе посвятив, дав тебе за пророка народам!
JER|1|6|А я відповів: О, Господи, Боже, таж я промовляти не вмію, бо я ще юнак!...
JER|1|7|Господь же мені відказав: Не кажи: Я юнак, бо ти підеш до всіх, куди тільки пошлю Я тебе, і скажеш усе, що тобі накажу.
JER|1|8|Не лякайсь перед ними, бо Я буду з тобою, щоб тебе рятувати, говорить Господь!
JER|1|9|І простяг Господь руку Свою, і доторкнувсь моїх уст та й до мене сказав: Ось Я дав в твої уста слова Мої!
JER|1|10|Дивись, Я сьогодні призначив тебе над народами й царствами, щоб виривати та бурити, і щоб губити та руйнувати, щоб будувати й насаджувати!
JER|1|11|І було мені слово Господнє, говорячи: Що ти бачиш, Єреміє? А я відказав: Я бачу мигдалеву галузку.
JER|1|12|І сказав мені Господь: Ти добре бачиш, бо Я пильную Свого слова, щоб справдилось воно.
JER|1|13|І було мені слово Господнє подруге таке: Що ти бачиш? А я відказав: Я бачу кипляче горня, а перед його звернений з півночі на південь.
JER|1|14|І сказав мені Господь: З півночі відкриється зло на всіх мешканців землі.
JER|1|15|Бо ось Я покличу всі родини царств на півночі, говорить Господь, і вони поприходять, і поставлять кожен свого трона при вході до єрусалимських брам, і навколо при всіх мурах його та при всіх юдиних містах.
JER|1|16|І буду судитися з ними за всю їхню безбожність, що вони покинули Мене, і кадили іншим богам, і вклонялись чинам своїх рук.
JER|1|17|А ти підпережеш стегна свої та й устанеш, і будеш говорити їм усе, що Я накажу тобі; не бійся перед ними, щоб Я не злякав тебе перед ними!
JER|1|18|Бо Я ось сьогодні поставив тебе містом твердинним, і залізним стовпом, і мідяними мурами проти всієї цієї землі, проти царів Юди, проти його князів, проти його священиків та проти народу цієї землі.
JER|1|19|І будуть вони воювати з тобою, та не переможуть тебе, бо Я із тобою, говорить Господь, щоб тебе рятувати!
JER|2|1|І було мені слово Господнє, говорячи:
JER|2|2|Іди, і проголоси до вух дочки Єрусалиму, говорячи: Так говорить Господь: Я згадав тобі ласку юнацтва твого, ту любов, коли ти наречена була та за Мною ходила в пустині, в землі незасіяній.
JER|2|3|Ізраїль то святість для Господа, початок врожаю Його. Всі, що їли його, завинили, зло прийде на них, говорить Господь.
JER|2|4|Послухайте слова Господнього, доме Яковів та всі роди дому Ізраїля!
JER|2|5|Так говорить Господь: яку кривду знайшли батьки ваші в Мені, що вони віддалились від Мене й пішли за марнотою, і стали марними?
JER|2|6|І не спитали вони: де Господь, що нас вивів із краю єгипетського, що провадив Він нас по пустині, по землі степовій, повній ям, по краю сухому та темному, по краю, що в ньому ніхто не ходив, і що там не осілась людина?
JER|2|7|І впровадив Я вас до родючого Краю, щоб їсти плоди його й добра його. І ви прибули й занечистили землю Мою, і зробили гидотою спадщину Мою...
JER|2|8|Священики не повіли: де Господь? А ті, хто тримає Закона, Мене не пізнали, і пастирі повідпадали від Мене, а пророки Ваалом пророкували, та за тими пішли, хто вам не допоможе...
JER|2|9|Тому то судитися буду ще з вами, говорить Господь, і з синами синів ваших буду судитись!
JER|2|10|Бо перейдіть острови хіттеян, і побачте, і до Кедару пошліть, та пригляньтеся добре й побачте, чи було там таке, як оце?
JER|2|11|Чи змінив люд богів, хоч не Бог вони? А народ Мій змінив свою славу на те, що не помагає!...
JER|2|12|Здивуйтеся цим, небеса, і затремтіть, і злякайтесь над міру, говорить Господь!
JER|2|13|Бо дві речі лихі Мій народ учинив: покинули Мене, джерело живої води, щоб собі подовбати водозбори, водозбори поламані, що води не тримають.
JER|2|14|Чи Ізраїль Мій раб? Чи він теж кріпак, народжений вдома? Чому ж здобиччю він?
JER|2|15|На нього ревуть левчуки, видають голос свій, і його Край обернули в пустиню, спалили міста його, так що немає мешканця...
JER|2|16|Також сини Мемфіса й Тахпенеса на черепі паслися в тебе.
JER|2|17|Чи ж зробило тобі це не те, що покинув ти Господа, Бога свого, що провадив тебе по дорозі?
JER|2|18|І тепер що тобі до дороги в Єгипет? Щоб пити воду з Шіхору? І що тобі до дороги в Ашшур? Щоб пити воду з Ріки?
JER|2|19|Хай карає тебе твоє зло, і відступства твої хай картають тебе, і пізнай та побач, що лихе та гірке це, що кинув ти Господа, Бога свого, і страху Мого над тобою нема, говорить Господь, Бог Саваот.
JER|2|20|Бо віддавна зламала ти, дочко Сіону, ярмо своє, пірвала свої поворозки й сказала: Не буду служити! Бо на кожному взгір'ї високому, і під кожним зеленим деревом ти клалась блудницею...
JER|2|21|А Я ж посадив був тебе виноградом добірним, увесь він насіння правдиве! І як ти змінилась Мені на виродка винограду чужого?
JER|2|22|Тому то хоч би ти й помилася лугом, і мила багато собі зажила б, проте плямою буде вина твоя перед обличчям Моїм, говорить Господь Бог!
JER|2|23|Як ти зможеш сказати: Я не стала нечистою, за Ваалами я не ходила? Подивись на дорогу свою, у долині, чого ти наробила, пустотлива верблюдко, що крутиш дороги свої!
JER|2|24|Ти як дика ослиця, яка до пустині привикла, що вітер втягає в жаданні своєї душі, хто заверне її в час її похотливости? Усі, хто шукає її, не помучаться, знайдуть її в її місяці!
JER|2|25|Стримуй ногу свою, щоб не бути їй босою, і від прагнення горло своє. А ти кажеш: Пропало, вже ні, бо я покохала чужих і за ними піду...
JER|2|26|Як для злодія сором, коли буде зловлений, так себе осоромив Ізраїлів дім, вони та царі їхні, їхні зверхники, й їхні священики, й їхні пророки,
JER|2|27|що говорять до дерева: Ти батько мій, а до каменя: Ти мене породив. Бо до Мене вони повернулись плечима, а не обличчям, а за час свого лиха говорять: Устань та спаси нас!
JER|2|28|А де ж твої боги, яких наробив ти собі? Хай устануть вони, якщо можуть спасти тебе в час твого лиха, бож в тебе богів, скільки міст твоїх, Юдо!
JER|2|29|Чого вам зо Мною змагатися? Усі ви відпали від Мене, говорить Господь.
JER|2|30|Надармо Я бив синів ваших, науки вони не взяли, а ваших пророків ваш меч поз'їдав, немов лев той винищувач!
JER|2|31|О ви, покоління, почуйте це слово Господнє: Чи пустинею був для Ізраїля Я? Чи може землею великої темряви? Чому ж каже народ Мій: Ми вільно буяємо, вже не прийдемо до Тебе?
JER|2|32|Чи панна забуде оздобу свою, наречена про стрічки свої? А народ Мій про Мене забув незчисленні вже дні!
JER|2|33|Як ти вправно дорогу свою повела, щоб шукати кохання! Тому то дороги свої призвичаїла ти до злочинства,
JER|2|34|і навіть на полах одежі твоєї знаходиться кров душ убогих невинних, яких не зловила на вчинку гарячому, але понад усім тим
JER|2|35|ти кажеш: Невинна я, Його гнів відвернувся від мене направду... Ось Я буду змагатись з тобою за те, що ти кажеш: Я не прогрішила!
JER|2|36|Нащо тиняєшся ти, і міняєш дорогу свою? Таж ти посоромлена будеш Єгиптом, як ти посоромлена від Асирії!
JER|2|37|І звідти ти вийдеш, заламуючи свої руки на своїй голові, бо повідкидав Господь тих, на кого ти надіялася, і не будеш ти мати в них успіху...
JER|3|1|І було мені слово Господнє, говорячи: Як відпустить хто жінку свою, й вона піде від нього, та стане за жінку для іншого чоловіка, чи вернеться ще він до неї? Чи ж не стане зовсім обезчещеною оця жінка? Ти ж перелюб чинила з коханцями багатьома, і тобі повертатись до Мене? говорить Господь.
JER|3|2|Зведи свої очі на гори порожні й дивися, де перелюбу ти не чинила? Ти для них по дорогах сиділа, немов той араб на пустині, і збезчестився край твоїм блудом та лихом твоїм!
JER|3|3|І дощі були стримувані, і не було дощу пізнього, проте мала ти чоло блудниці, і стратила сором...
JER|3|4|Чи ж кликати віднині не будеш до Мене: Отче мій, Ти юнацтва мого Провідник!
JER|3|5|Чи Він пам'ятатиме вічно про гнів, чи назавжди його стерегтиме? Таке ти говориш, і безмежно зло чиниш...
JER|3|6|І сказав до мене Господь за днів царя Йосії: Чи ти бачив, що зробила невірна дочка Ізраїлева? Вона ходила на кожну високу гору, і під кожне зелене дерево, і блудодіяла там...
JER|3|7|Я думав: Як зробить вона все оце, то до Мене повернеться; та вона не вернулась, і бачила це сестра її зрадниця, Юдея.
JER|3|8|І побачила Юдея, що за все те, що перелюб чинила невірна дочка Ізраїлева, відпустив Я її, і дав їй листа розводового. Та зрадлива сестра її, дочка Юдина, не побоялася й пішла, і блудливою стала й вона...
JER|3|9|І сталось від розголосу про перелюб її, збезчестила вона землю, і перелюб чинила з камінням та з деревом.
JER|3|10|І також при всьому цьому не вернулась до Мене зрадлива сестра її, дочка Юди, усім своїм серцем, а тільки вдавала, говорить Господь...
JER|3|11|І промовив до мене Господь: Невірна дочка Ізраїлева всправедливила душу свою більш від зрадливої дочки Юди.
JER|3|12|Піди, і проголосиш слова ці на північ та й скажеш: Вернися, відступна дочко Ізраїлева! говорить Господь. Не зверну Я Свого обличчя у гніві на вас, бо Я милостивий, говорить Господь, і не буду повік стерегти Свого гніву.
JER|3|13|Тільки пізнай же провину свою, бо ти проти Господа, Бога свого повстала, і грішила з чужими під деревом кожним зеленим, і Мого голосу ви не почули, говорить Господь.
JER|3|14|Верніться, діти невірні, говорить Господь, бо Я вам Господар, та візьму вас по одному з міста, а з роду по два, і вас поведу до Сіону!
JER|3|15|І дам пастирів вам згідно з серцем Своїм, і вони будуть пасти вас умінням та розумом.
JER|3|16|І буде, коли ви розмножитеся та розплодитеся на землі за цих днів, говорить Господь, не скажуть уже: ковчег заповіту Господнього, і він вже не прийде на серце, і його пам'ятати не будуть, і більше не буде він зроблений...
JER|3|17|Того часу назвуть Єрусалима: Господній престол, і до нього, до Єрусалиму згромаджені будуть народи усі ради Ймення Господнього, і більше не підуть вони за впертістю серця лихого свого...
JER|3|18|Тими днями дім Юдин із домом Ізраїля підуть і разом прибудуть з північного краю до краю, що вашим батькам на спадок Я дав.
JER|3|19|І Я був подумав: як поставлю тебе Я посеред синів і дам тобі край пожаданий, найкращу спадщину народів? І Я думав: ви будете звати Мене: Мій Отче, і не відвернетеся ви від Мене.
JER|3|20|Справді, як зраджує жінка свого чоловіка, так ви Мене зрадили, доме Ізраїлів! каже Господь.
JER|3|21|Чути голос на лисих горах, плач благальний синів Ізраїлевих, вони бо скривили дорогу свою, забули про Господа, Бога свого:
JER|3|22|Верніться, невірні сини, усі ваші відступства Я вилікую! Ось прийшли ми до Тебе, бо Ти Господь, Бог наш!
JER|3|23|Справді, неправда ті пагірки, той гомін на горах, справді, в Господі, Богові нашім, спасіння Ізраїлеве!
JER|3|24|А той сором пожер працю наших батьків від нашої молодости, їхню худобу дрібну й їхню худобу велику, синів їхніх та їхніх дочок.
JER|3|25|Лежимо ми у соромі нашому, і нас покриває ця наша неслава, бо ми прогрішилися Господу, Богові нашому, ми й батьки наші, від нашої молодости й до сьогодні, і не слухали голосу Господа, нашого Бога!...
JER|4|1|Якщо ти, Ізраїлю, вернешся, каже Господь, до Мене ти вернешся, і якщо ти відкинеш із-перед обличчя Мого гидоти свої, то не будеш тинятись!
JER|4|2|І якщо ти присягнеш Як живий Господь правдою й правом та справедливістю, то будуть Ним благословлятись народи, і хвалитись Ним будуть.
JER|4|3|Бо так каже Господь мужам Юди та Єрусалиму: Оріть собі на цілині, і не сійте в тернину!
JER|4|4|Обрізуйтеся Господеві, й усуньте із ваших сердець крайні плоті, юдеї та мешканці Єрусалиму, щоб не вийшла, немов той огонь, Моя лютість, і буде палати вона, і не буде кому погасити через злі ваші вчинки!
JER|4|5|Оповістіте в Юдеї та в Єрусалимі звістіть та й скажіть: Засурміте в сурму у краю! Кричіть гучним голосом та говоріть: Зберіться та підемо до міст до твердинних!
JER|4|6|Підійміте прапор до Сіону, поспішайте, не станьте, бо з півночі зло приведу, і велике нещастя...
JER|4|7|Лев виходить із своєї гущавини, і той, хто нищить народи, вирушає із місця свого, щоб твій край обернути на руїну, і спустошені будуть міста твої, так що забракне і мешканця!...
JER|4|8|Отож, опережіться веретами, плачте та голосіть, бо лютість Господнього гніву від нас не відвернеться!
JER|4|9|І станеться в день той, говорить Господь, згине розум царя і розум князів, і остовпіють священики, а пророки здивуються
JER|4|10|й скажуть: О Господи, Боже, справді обманений сильно народ цей та Єрусалим, коли казано: Буде вам мир, а меч доторкнувся ось аж до душі!...
JER|4|11|Того часу народові цьому та Єрусалимові сказане буде: Ось вітер палкий з лисих гір на пустині, на дорозі дочки Мого люду, не на віяння й не на очищення він!
JER|4|12|Та вітер сильніший від цього прибуде Мені, і над ними Я суд прокажу...
JER|4|13|Ось він прийде, як хмари, й як буря його колесниці, від орлів швидші коні його: Горе нам, бо спустошені будемо ми!...
JER|4|14|Обмий серце своє від лихого, о Єрусалиме, щоб був ти врятований! Аж доки в тобі пробуватимуть думки марноти твоєї?
JER|4|15|Бо голос доносить із Дану й звіщає погибіль з Єфремових гір...
JER|4|16|Пригадайте народам оце, сповістіть ось про Єрусалим: Приходять з далекого краю його облягати, і здіймають свій крик на юдейські міста!
JER|4|17|Як сторожа полів, навколо оточать його, бо він Мені був неслухняний, говорить Господь!
JER|4|18|Дорога твоя й твої вчинки тобі це зробили, це лихо твоє: бо гірке, бо торкнуло воно аж до серця твого...
JER|4|19|Ой, утробо моя, ти утробо моя, я тремчу! Біль серце стискає мені, і трепоче мені моє серце!... Не можу мовчати, бо вчула душа моя голос сурми, гук війни!
JER|4|20|Біда на біду прикликається, вся бо земля поруйнована буде, спустошені будуть зненацька намети мої, вмить завіси мої...
JER|4|21|Аж доки я бачити прапора буду, буду чути голос сурми?
JER|4|22|Тому, що народ мій безглуздий, він не знає Мене: вони нерозумні сини й нерозважні вони, мудрі вони, щоб чинити лихе, та не вміють чинити добра!
JER|4|23|Дивлюся на землю, аж ось порожнеча та пустка, і на небо й нема його світла!
JER|4|24|Дивлюся на гори, аж ось вони трусяться, і всі згір'я хитаються!
JER|4|25|Дивлюся, аж ось вже немає людини, і порозліталось все птаство небесне.
JER|4|26|Дивлюся, аж ось край родючий пустинею став, а міста його знищені всі від обличчя Господнього, від полум'я гніву Його...
JER|4|27|Бо Господь так прорік: Спустошенням стане ввесь край, та кінця йому ще не вчиню!
JER|4|28|І буде в жалобі земля через це, і затьмариться небо вгорі, бо Я говорив, що задумав, і не пожалую, і не відступлюся від того...
JER|4|29|Від гуркотнечі їздця та стрільця побіжить усе місто, повтікають в гущавини й злізуть на скелі... Всі міста покинуті, і немає нікого, хто мешкав би в них...
JER|4|30|А ти, поруйнована, дочко Сіону, що будеш робити? Хоч ти зодягаєш себе в кармазин, хоч прикрашуєшся золотою оздобою, хоч очі свої підмальовуєш фарбою, та надаремно прикрашуєшся: обридили тобою коханці твої, на життя твоє важать вони!
JER|4|31|Бо чую Я крик, немов породіллі, чую стогін, мов первістки, голос Сіонської дочки, вона стогне, заломлює руки свої та голосить: Ой, горе мені, бо попало життя моє вбивникам!...
JER|5|1|Помандруйте по вулицях Єрусалиму, і розгляньтеся та розпізнайте, і на майданах його пошукайте: чи не знайдете там людини, чи нема там такого, що чинить за правом, що правди шукає, то Я їм пробачу!
JER|5|2|Коли ж вони кажуть: Як живий Господь, то справді клянуться неправдою.
JER|5|3|Хіба ж очі Твої не для правди, о Господи? Уразив Ти їх, але їм не болить, понищив Ти їх, та відмовились узяти поуку вони, обличчя свої поробили від скелі твердішими, відмовилися навернутись!
JER|5|4|А Я думав: Це прості лиш люди, безглузді, вони бо не знають дороги Господньої, права Бога свого.
JER|5|5|Піду но собі до вельможних і з ними помовлю, бо знають дорогу Господню вони, право Бога свого, та й вони усі разом зламали ярмо, а шлеї пірвали!
JER|5|6|Тому лев лісовий їх поб'є, погубить їх вовк степовий, пантера чигає на їхні міста: кожен, хто вийде із них, пошматований буде, бо помножились їхні гріхи, їхні відступства численними стали!
JER|5|7|Хіба через це Я пробачу тобі: твої діти Мене полишили, і присягаються тим, хто не Бог. Я їх нагодував, а вони чужоложать і натовпом ходять до дому блудниці,
JER|5|8|волочаться, мов жеребці відгодовані: кожен ірже до жони свого ближнього...
JER|5|9|Чи ж оцього Я не покараю? говорить Господь. І хіба над народом, як цей, не помститься душа Моя?
JER|5|10|Зберіться на мури його та й понищте, але не вчиняйте кінця їм! Усуньте підпори його, бо вони не для Господа,
JER|5|11|бо зраджуючи, Мене зрадив Ізраїлів дім та дім Юдин, говорить Господь.
JER|5|12|Вони відцуралися Господа та говорили: Немає Його, й зло не прийде на нас, ні меча, ані голоду ми не побачимо!
JER|5|13|А пророки поробляться вітром, і немає в них слова Господнього, отак їм пороблено буде!
JER|5|14|Тому вирікає отак Господь Бог Саваот: За те, що говорите слово таке, ось Я в уста твої вкладу слово Своє за огонь, а народ цей то дрова, і він пожере їх!
JER|5|15|Ось Я приведу іздалека народа на вас, о доме Ізраїлів, каже Господь, це сильний народ, стародавній це люд, люд, що мови його ти не знаєш, і не зрозумієш, що він говоритиме.
JER|5|16|Його сагайдак, як відчинений гріб, усі хоробрі вони.
JER|5|17|І він пожере твоє жниво та хліб твій, поїсть він синів твоїх та дочок твоїх, худобу дрібну та худобу велику твою пожере, з'їсть твого виноградника й фіґу твою, понищить мечем твердинні міста твої, на які ти надієшся...
JER|5|18|Та й за тих днів, говорить Господь, не зроблю Я із вами кінця!
JER|5|19|І буде, як скажуть: За що Господь, Бог наш зробив нам усе це? то ти скажеш до них: Як Мене ви покинули, і служите в вашому краї богам чужоземним, так чужинцям служити ви будете в краї не вашому!...
JER|5|20|Сповістіть в домі Якова це, та оголосіть це в Юдеї, говорить Господь.
JER|5|21|Почуй же оце, ти народе безумний й безсердий, який має очі й не бачить, має вуха й не чує!
JER|5|22|Чи Мене ви боятись не будете, каже Господь, чи тремтіти не будете перед лицем Моїм? Мене, що пісок поклав за границю для моря, за вічну межу, якої воно не перейде: хоч повстануть, та не переможуть, і шумітимуть хвилі його, але не переступлять її!
JER|5|23|А серце в народа цього неслухняне та непокірне, відпали вони та й пішли.
JER|5|24|І не сказали вони в своїм серці: Біймося ж Господа, нашого Бога, який дає дощ, дощ ранній та пізній часу його, стереже нам уставлені тижні для жнив.
JER|5|25|Ваші провини оце відхилили, а ваші гріхи від вас стримали цеє добро.
JER|5|26|Бо в народі Моєму безбожники є, чигають вони, немов той птахолов, вони сітки розставили, хапають людей...
JER|5|27|Як клітка, наповнена птахами, так доми їхні повні омани, тому повиростали та збагатились вони!
JER|5|28|Потовстіли вони та погладшали, переступають також міру злого, справедливо вони не судили сирітського суду, і мають поводження! і не помагають убогим у їхній справі.
JER|5|29|Чи ж оцього Я не покараю? говорить Господь. І хіба над народом, як цей, не помститься душа Моя?
JER|5|30|Чудне та страшне стало в краї:
JER|5|31|пророки віщують неправду, при помочі їхній панують священики, і народ Мій оце так кохає! І що зробите ви, як кінець тому прийде?
JER|6|1|Утікайте, сини Веніямина, з середини Єрусалиму, і засурміте в сурму у Текої, і знак підійміть на Бет-Гаккерем, бо з півночі грізно підноситься зло та велике нещастя!
JER|6|2|І викореню Я Сіонську дочку, вродливу та випещену.
JER|6|3|Пастухи поприходять до неї з своїми стадами, понапинають намети навколо при ній, кожен місце своє випасатиме.
JER|6|4|Приготуйте війну проти неї, вставайте та вдармо опівдні! Горе нам, бо минає вже день, бо вже тягнуться тіні вечірні!
JER|6|5|Уставайте та підемо вночі і понищмо палати її!
JER|6|6|Бо так промовляє Господь Саваот: Постинайте дерева та вала насипте при Єрусалимі! Він те місто, що має зруйноване бути, в ньому повно насильства:
JER|6|7|як виприскує воду свою джерело, так виприскує він своє зло... Насилля й грабіж чуті в ньому, перед обличчям Моїм безперестань хвороба та рана...
JER|6|8|Будь навчений, Єрусалиме, щоб душа Моя не відвернулась від тебе, щоб тебе не вчинив Я спустошенням, незаселеним краєм!
JER|6|9|Так говорить Господь Саваот: Позбирають дорешти останки Ізраїля, мов виноградові рештки, простягни свою руку, немов виноградар по грона!
JER|6|10|До кого я буду казати та свідчити буду, і слухатимуть? Необрізане ось їхнє вухо і слухати уважно не можуть вони, ось слово Господнє для них стало посміхом вони не жадають його!
JER|6|11|І гніву Господнього повен я став, змучився я, його стримуючи, на вулиці виллю його на дітей та на збір юнаків одночасно, бо схоплені будуть чоловік із жінкою, старий із віджилим літа,
JER|6|12|і дістануться іншим доми їхні, теж поля та жінки... Бо Я руку Свою простягну на мешканців цієї землі, говорить Господь.
JER|6|13|Бо вони від малого свого й до великого, усі пожадливі на зиски, і від пророка та аж до священика роблять неправду...
JER|6|14|І рани народу Мого легковажно лікують, говорячи: Мир, мир, а миру нема!
JER|6|15|Чи вони засоромилися, що гидоту робили? не засоромилися ані трохи вони й застидатись не вміють... Тому то впадуть між упалими в часі, коли їх навіщу Я, спіткнуться, говорить Господь.
JER|6|16|Так говорить Господь: На дорогах спиніться та гляньте, і спитайте про давні стежки, де то добра дорога, то нею ідіть, і знайдете мир для своєї душі! Та вони відказали: Не підемо!
JER|6|17|І Я сторожів був поставив над вами, говорячи: Прислухайтесь до голосу сурми! Та вони відказали: Не будем прислухуватись!
JER|6|18|Тому слухайте, люди, і пізнай, ти громадо, що станеться з ними.
JER|6|19|Послухай, ти земле: Ось Я веду на народ цей лихе, плід їхніх думок, бо до слів Моїх не прислухались вони, а Законом Моїм погордили!
JER|6|20|Навіщо Мені те кадило, що з Шеви приходить, запашний очерет із далекого краю? Цілопалення ваші не любі Мені, ваші ж жертви Мені не приємні!
JER|6|21|Тому то Господь каже так: Ось Я дам спотикання оцьому народові, і спіткнуться об них разом ваші батьки та сини, сусід та приятель його, і загинуть!
JER|6|22|Так говорить Господь: Ось приходить народ із північного краю, і збуджується люд великий із кінців землі.
JER|6|23|Лука та ратище міцно тримають, жорстокі вони й милосердя не мають, їхній голос, як море реве, і гарцюють на конях вони... Ушикований, мов чоловік той до бою, на тебе, о дочко Сіону!
JER|6|24|Як почули ми звістку про нього, омліли нам руки, обняла нас тривога та біль, немов в породіллі...
JER|6|25|Не виходьте на поле й не йдіте дорогою, бо в ворога меч та страхіття навколо!
JER|6|26|Дочко народу Мого, веретою підпережись та качайся у попелі! Справ жалобу собі, немов над однородженим, голосіння гірке, бо прийде зненацька руїнник на нас!
JER|6|27|Я дав був тебе випробовувачем у народі Моїм, за твердиню, щоб ти знав і випробовував їхню дорогу.
JER|6|28|Вони всі відступники над відступниками, чинять наклепи, усі вони мідь та залізо, вони згубники!...
JER|6|29|Спалилося духало, від огню зникло оливо, надармо старанно розтоплювано, бо злих не відділено...
JER|6|30|Сріблом відкиненим названо їх, бо Господь їх відкинув.
JER|7|1|Слово, що було до Єремії від Господа, говорячи:
JER|7|2|Стань у брамі Господнього дому, і прокажеш там слово оце та промовиш: Послухайте слово Господнє, ввесь Юдо, що ходите брамами цими вклонятися Господу.
JER|7|3|Так говорить Господь Саваот, Бог Ізраїлів: Поправте дороги свої й свої вчинки, й Я зроблю, що ви житимете на цім місці!
JER|7|4|Не надійтесь собі на слова неправдиві, щоб казати: Храм Господній, храм Господній, храм Господній отут!
JER|7|5|Бо якщо ви насправді поправите ваші дороги та ваші діла, якщо один одному будете справді чинити справедливо,
JER|7|6|не будете тиснути чужинця, сироту та вдову, не будете лити невинної крови на місці цьому, і за іншими богами вслід не підете собі на біду,
JER|7|7|то зроблю, що ви пробуватимете на цім місці, у Краю, що його дав Я вашим батькам відвіку навіки!
JER|7|8|Ось собі ви надієтеся на слова неправдиві, які не допоможуть:
JER|7|9|Чи ви будете красти, вбивати й перелюб чинити, і присягати фальшиво, й кадити Ваалові, і ходити за іншими богами, яких ви не знаєте,
JER|7|10|а потім ви прийдете й станете перед обличчям Моїм у цім домі, що зветься Ім'ям Моїм, і скажете: Урятовані ми, щоб чинити гидоти всі ці?
JER|7|11|Чи вертепом розбійників став оцей дім, що Ім'я Моє кличеться в ньому, на ваших очах? І Я оце бачу, говорить Господь...
JER|7|12|Бо підіть но до місця Мого, що в Шіло, де Я спочатку вчинив був перебування для Ймення Свого, і побачите, що вчинив Я йому через лукавство Мого народу Ізраїлевого...
JER|7|13|Тепер же за те, що ви робите всі оці вчинки, говорить Господь, і що Я говорив був до вас, промовляючи пильно, але ви не слухали, і кликав Я вас, та ви не відказали,
JER|7|14|то зроблю цьому домові, що кликалось в ньому Ім'я Моє, що на нього надієтесь ви, і місцю цьому, що Я дав його вам та вашим батькам, так само, як Я був зробив для Шіло,
JER|7|15|і відкину Я вас від обличчя Свого, як відкинув усіх ваших братів, усе насіння Єфремове!...
JER|7|16|А ти не молись за народ цей, і благання й молитви за них не здіймай, і Мене не проси, бо не вислухаю Я тебе!
JER|7|17|Хіба ти не бачиш, що роблять вони в містах Юдиних та на вулицях Єрусалиму:
JER|7|18|Діти дрова збирають, а батьки розкладають огонь, жінки ж місять тісто, щоб спекти калачів тих жертовних небесній цариці, і ллють литі жертви для інших богів, на досаду Мені...
JER|7|19|Та хіба ображають Мене, говорить Господь? Хіба не себе самих, щоб сором покрив їхні обличчя?
JER|7|20|Тому Господь Бог промовляє отак: Ось ллється Мій гнів і Моя лють на це місце, на людину й худобу, і на польові дерева та на земні плоди, і палатиме він, і не згасне!
JER|7|21|Так говорить Господь Саваот, Бог Ізраїлів: Додайте свої цілопалення до жертов ваших, і їжте м'ясо,
JER|7|22|бо Я не говорив батькам вашим, і не наказував їм того дня, як виводив їх із краю єгипетського, про справи цілопалення й жертви.
JER|7|23|Бо лиш справу оцю Я звелів їм, говорячи: Слухайтеся Мого голосу, і Я буду вам Богом, а ви будете народом Моїм, і ходіть усією дорогою, про яку накажу вам, щоб вам було добре.
JER|7|24|Та не слухали й не нахилили вони свого вуха, а ходили за радами та за упертістю серця лихого свого, і стали до Мене плечима, а не обличчям.
JER|7|25|Від того дня, коли ваші батьки вийшли з краю єгипетського, аж до дня цього, посилав Я до вас усіх Своїх рабів пророків, посилав щодня пильно.
JER|7|26|Та вони не слухалися Мене, і вуха свого не схиляли, і показали себе твердошийними, зло чинили ще більш від батьків своїх...
JER|7|27|І ти будеш казати їм ці всі слова, та не будуть вони тебе слухати, і будеш ти кликати до них, та вони тобі відповіді не дадуть...
JER|7|28|І скажеш до них: Оце той народ, що не слухався голосу Господа, Бога свого, і поуки не брав, загинула правда, і зникла з їхніх уст...
JER|7|29|Обстрижи ти волосся своє та й відкинь, на лисих горах здійми жалісний спів, бо відкинув Господь і покинув плем'я Свого гніву!
JER|7|30|Бо Юдині сини чинять зло в Моїх очах, говорить Господь, поклали гидоти свої в тому домі, що в нім кликалося Моє Ймення, щоб збезчестити його...
JER|7|31|І побудували ті жертовні пагірки Тофета, що в долині Бен-Гіннома, щоб палити синів своїх та дочок своїх на огні, чого Я не наказував, і що на серце Мені не приходило...
JER|7|32|Тому то приходять ось дні, говорить Господь, що не буде вже кликатись Тофет місце це чи Долина Бен-Гіннома, а тільки Долина вбивства, і будуть ховати у Тофеті через брак місця на погреб.
JER|7|33|І стане труп цього народу за стерво небесному птаству та земній звірині, і не буде, хто б їх відстрашив!...
JER|7|34|І спиню в містах Юдиних та на вулицях Єрусалиму голос радісний і голос веселий, голос молодого та голос молодої, бо руїною стане цей Край!
JER|8|1|Того часу, говорить Господь, повитягують кості царів Юди та кості його князів, і кості священиків, і кості пророків, і кості мешканців Єрусалиму з їхніх гробів,
JER|8|2|і порозкладають їх перед сонцем і перед місяцем, та перед усіма небесними світилами, яких вони кохали та служили їм, і що йшли за ними, і що зверталися до них, і що вклонялися їм. Не будуть вони зібрані й не будуть поховані, гноєм стануть вони на поверхні землі!
JER|8|3|І смерть буде ліпша від життя для всієї решти позосталих зо злого цього роду, по всіх цих місцях позосталих, куди Я їх повиганяв, говорить Господь Саваот.
JER|8|4|І скажеш до них: Так говорить Господь: Хіба падають і не встають? Хіба хто відступить, то вже не вертається?
JER|8|5|Чому відступив оцей єрусалимський народ усевічним відступленням? Міцно схопились вони за оману, не хочуть навернутись.
JER|8|6|Прислухався Я й слухав: неправду говорять, немає нікого, хто б каявсь у своєму лукавстві, говорячи: Що я зробив? Кожен з них обертається до свого бігу, мов той кінь, що женеться у бій...
JER|8|7|І відає бусел у повітрі умовлений час свій, а горлиця й ластівка та журавель стережуть час прилету свого, а народ Мій не знає Господнього права!...
JER|8|8|Як ви скажете: Ми мудреці, і з нами Господній Закон? Ось справді брехнею вчинило його брехливе писарське писальце!
JER|8|9|Засоромлені ці мудреці, збентежилися й були схоплені. Ось вони слово Господнє відкинули, що ж за мудрість ще мають вони?
JER|8|10|Тому їхніх жінок віддам іншим, а їхні поля здобувцям, бо вони від малого та аж до великого усі віддались користолюбству, від пророка та аж до священика чинять неправду!...
JER|8|11|І легенько лікують нещастя народу Мого, говорячи: Мир, мир, а миру нема!
JER|8|12|Чи вони засоромилися, що гидоту робили? Ні трохи вони не засоромилися, і застидатись не вміють, тому то впадуть між упалими в часі навіщення їх, спіткнуться, говорить Господь...
JER|8|13|Зберу їх дощенту, говорить Господь: не буде ягід у них на винограді, і не буде на фіґовім дереві фіґ, а їхнє листя пов'яне, і пошлю їм таких, що їх поїдять...
JER|8|14|Пощо ми сидимо? Збирайтесь та підемо в твердинні міста та й погинемо там, бо Господь, Бог наш, учинив, що ми згинемо, і напоїв нас водою трійливою, бо ми Господеві згрішили...
JER|8|15|Ми миру чекали, й немає добра, часу вилікування й ось жах!
JER|8|16|Чути фиркання коней його аж від Дану, від гуку іржання його жеребців уся земля затремтіла! І прийдуть вони, й пожеруть усю землю та повню її, місто й тих, хто замешкує в ньому...
JER|8|17|Бо ось Я пошлю проти вас тих вужів та гадюк, що немає закляття на них, і вони вас кусатимуть, каже Господь!
JER|8|18|Яка моя втіха у смутку? Болить мені серце моє...
JER|8|19|Ось голосіння дочки Мого народу з далекого краю: Чи Господь не в Сіоні? Чи не в нім його Цар? Нащо Мене розгнівили своїми бовванами, тими чужими марнотами?
JER|8|20|Минули жнива, покінчилося літо, а ми не спасені...
JER|8|21|Через нещастя дочки народу мого знещасливлений я, і міцно страхіття мене обняло...
JER|8|22|Чи немає бальзаму в Ґілеаді? Чи ж немає там лікаря? Чому нема вилікування для доньки народу Мого?
JER|9|1|(8-23) Ой, коли б голова моя стала водою, а око моє за джерело сльози, то я плакав би вдень та вночі над побитими доньки народу мого!...
JER|9|2|(9-1) Ой, коли б на пустині нічліг подорожніх я мав, тоді б я покинув народа свого, і пішов би від них, бо вони перелюбники всі, збори зрадників!
JER|9|3|(9-2) Вони напинають свого язика, немов лука свого, для неправди, міцніють вони на землі не для правди, бо від злого до злого ідуть і не знають Мене, говорить Господь!
JER|9|4|(9-3) Один одного остерігайтесь, і не покладайтесь на жодного брата, кожен бо брат обманити обманить, і приятель кожен обмовник!
JER|9|5|(9-4) Один одного зводить, і правди не кажуть, привчили свого язика говорити неправду, помучилися, лихо чинячи!
JER|9|6|(9-5) Серед омани твоє проживання, через оману не хочуть пізнати Мене, говорить Господь.
JER|9|7|(9-6) Тому так промовляє Господь Саваот: Ось Я їх перетоплюю та випробовую їх, бо що маю вчинити Я ради дочки Свого люду?
JER|9|8|(9-7) Їхній язик смертоносна стріла, він оману говорить: устами своїми говорить із ближнім про мир, а в нутрі своєму кладе свою засідку...
JER|9|9|(9-8) Чи ж за це Я їх не покараю? говорить Господь. Хіба ж над народом, як цей, непомститься душа Моя?
JER|9|10|(9-9) Я плач та ридання здійму над оцими горами, і спів жалобний понад степовими лугами, вони бо попалені так, що ними не ходить ніхто, і реву худоби не чути: від птаства небесного й аж до худоби розбіглося все, відійшло!
JER|9|11|(9-10) І Я Єрусалим на руїни віддам, на мешкання шакалів, а юдські міста на спустошення дам, і не буде мешканця у них!
JER|9|12|(9-11) Хто муж мудрий, який зрозумів би оце, і до кого Господні уста промовляли, щоб вияснить те, за що згинув цей Край, за що спалений він, як пустиня, і що нею не ходить ніхто?
JER|9|13|(9-12) А Господь відказав: За те, що вони покинули Закона Мого, що Я дав перед ними, і не слухалися Мого голосу, і не ходили за ним, за Законом,
JER|9|14|(9-13) а ходили за впертістю серця свого й за Ваалами, що навчили про них їхні батьки...
JER|9|15|(9-14) Тому так промовляє Господь Саваот, Бог Ізраїлів: Ось Я їх, цей народ, полином нагодую й водою отруйною їх напою!
JER|9|16|(9-15) І розпорошу Я їх серед народів, яких ні вони, ні батьки їхні не знали, і пошлю Я за ними меча, аж поки не вигублю їх!
JER|9|17|(9-16) Так говорить Господь Саваот: Розгляньтеся та голосільниць покличте, і нехай вони прийдуть, і пошліте до мудрих жінок, і вони поприходять!
JER|9|18|(9-17) І хай поспішають, і хай спів жалоби над ними підіймуть, і хай наші очі зайдуться сльозою, а з наших повіків вода хай тече!
JER|9|19|(9-18) Бо почується голос жалобного співу з Сіону: Як ми попустошені, як посоромлені дуже!... Бо ми покинули свій край, бо покинули місце свого пробування...
JER|9|20|(9-19) Тож почуйте, жінки, слово Господа, і хай ваше ухо візьме слово уст Його, і навчіть дочок ваших жалобного співу, й одна одну жалобної пісні!
JER|9|21|(9-20) Бо смерть увійшла в наші вікна, до наших палат увійшла, щоб вирізати дітей з вулиці, із площ юнаків...
JER|9|22|(9-21) Кажи так: Говорить Господь: І нападає людського трупа, мов гною на полі, і мов тих снопів за женцем, і не буде кому позбирати!...
JER|9|23|(9-22) Так говорить Господь: Хай не хвалиться мудрий своєю премудрістю, і хай не хвалиться лицар своєю хоробрістю, багатий багатством своїм хай не хвалиться!
JER|9|24|(9-23) Бо хто буде хвалитись, хай хвалиться тільки оцим: що він розуміє та знає Мене, що Я то Господь, Який на землі чинить милість, правосуддя та правду, бо в цьому Моє уподобання, каже Господь!
JER|9|25|(9-24) Ось дні наступають, говорить Господь, і Я навіщу всіх обрізаних та необрізаних,
JER|9|26|(9-25) Єгипет та Юду, й Едома та Аммонових синів, і Моава та всіх, хто волосся довкола стриже, хто сидить на пустині, бо всі оці люди необрізані, а ввесь дім Ізраїлів необрізаносердий!...
JER|10|1|Послухайте слова того, що вам каже Господь, о доме Ізраїлів!
JER|10|2|Так говорить Господь: Не навчайтесь доріг цих народів, і небесних ознак не лякайтесь, бо тільки погани лякаються їх!
JER|10|3|Бо устави народів марнота вони, божок бо це дерево, з лісу вирубане, і це діло рук майстра сокирою!
JER|10|4|Сріблом та злотом його прикрашають, цвяхами та молотками прикріплюють їх, і він не захитається.
JER|10|5|Вони, як опудало на огірковім городі, й безмовні, і конче їх носять, бо не ходять вони. Не бійтеся їх, бо не вчинять лихого, і також учинити добро це не в їхній силі!
JER|10|6|Такого, як Ти, нема, Господи: Ти великий й велике Ім'я Твоє могутністю!
JER|10|7|Хто не буде боятись Тебе, Царю народів? Бо Тобі це належить, бо між усіма мудрецями народів і в усьому їхньому царстві немає такого, як Ти!
JER|10|8|Вони стали всі разом безумні й безглузді, наука марна оце дерево!
JER|10|9|Срібна бляха з Таршішу привезена, злото ж з Офіру, праця майстра й руки золотарської, блакить та пурпура їхня одіж, усі вони праця мистців.
JER|10|10|А Господь Бог правдивий, Він Бог Живий та Цар вічний! Від гніву Його затрясеться земля, і не знесуть Його гніву народи.
JER|10|11|Отак їм скажіть: боги, що неба й землі не вчинили, погинуть з землі та з-під неба цього!
JER|10|12|Своєю Він силою землю вчинив, Своєю премудрістю міцно поставив вселенну, і небо напнув Своїм розумом.
JER|10|13|Як голос Його забринить, у небесах шумлять води, а коли підіймає Він хмари із краю землі, коли блискавки чинить дощем та вітер виводить з криївок Своїх,
JER|10|14|тоді кожна людина дуріє в своєму знанні, усяк золотар посоромлений через боввана, бо відлив його це неправда, і немає в них духа!...
JER|10|15|Марнота вони, вони праця на сміх, в час навіщення їх вони згинуть!
JER|10|16|Не така, як оці, частка Яковова, бо Він все вформував, а Ізраїль племено спадку Його, Господь Саваот Його Ймення!
JER|10|17|Забери із землі свій товар, ти, що сидиш ув облозі!
JER|10|18|Бо Господь каже так: Ось цим разом Я кину мешканців цієї землі, мов із пращі, і притисну їх так, щоб пізнання знайшли...
JER|10|19|Ой, горе мені з-за нещастя мого, моя рана болюча! А я говорив: це хвороба моя, і знесу я її.
JER|10|20|Намета мого попустошено і зірвані всі мої шнури. Розійшлись мої діти від мене й нема їх, нема вже кому розтягнути намета мого та повісити завіси мої...
JER|10|21|Бо пастирі стали безглузді, і вони не звертались до Господа, тому не щастилося їм, і розпорошене все їхнє стадо...
JER|10|22|Голос звістки: Іде ось, і гуркіт великий з північного краю, щоб юдські міста обернути в спустошення, на мешкання шакалів...
JER|10|23|Знаю, Господи, я, що не в волі людини дороги її, не в силі людини, коли вона ходить, кермувати своїм кроком.
JER|10|24|Карай мене, Господи, тільки ж за судом, не гнівом Своїм, щоб не знищити мене!
JER|10|25|Вилий лютість Свою на народи, що не знають Тебе, та на роди, що Ймення Твого не кликали, що Якова з'їли й пожерли його, і погубили його, а мешкання його опустошили!...
JER|11|1|Слово, що було до Єремії від Господа, кажучи:
JER|11|2|Послухайте слів заповіту оцього, і будете їх говорити юдеям і мешканцям Єрусалиму,
JER|11|3|і скажеш ти їм: Так говорить Господь, Бог Ізраїлів: Проклята та людина, що не слухає слів заповіту цього,
JER|11|4|що його наказав був Я вашим батькам того дня, коли їх виводив із краю єгипетського, із залізного горна, говорячи: Слухайтеся Мого голосу, і робіть усе те, що Я накажу вам, і будете ви народом Моїм, а Я буду вам Богом,
JER|11|5|щоб Я виповнив присягу ту, якою Я вашим батькам присягав дати їм Край, що тече молоком, як сьогодні! А я відповів та сказав: Амінь, Господи!
JER|11|6|І промовив до мене Господь: Виголошуй оці всі слова по юдейських містах та на вулицях Єрусалиму, говорячи: Слухайтесь слів заповіту цього, і виконуйте їх!
JER|11|7|Бо направду засвідчив Я вашим батькам того дня, як виводив їх з краю єгипетського, і до сьогодні Я пильно засвідчую, кажучи: Слухайтеся Мого голосу!
JER|11|8|Та не слухали й не прихиляли вони свого вуха, і кожен ходив за упертістю злісного серця свого... І Я спровадив на них усі слова заповіту цього, що Я наказав був робити, вони ж не робили.
JER|11|9|І промовив до мене Господь: Знайдений бунт між юдеями та між мешканцями Єрусалиму!
JER|11|10|Повернулись вони до гріхів своїх давніх батьків, що слухатися Моїх слів не хотіли, і пішли за богами чужими, щоб їм служити. Дім Ізраїлів і дім Юдин зламали Мого заповіта, якого Я склав з їхніми батьками.
JER|11|11|Тому так промовляє Господь: Ось Я лихо на них наведу, що вийти із нього не зможуть, і кликати будуть до Мене, але не почую Я їх!
JER|11|12|І підуть юдейські міста та єрусалимські мешканці, і будуть кричати до богів, що їм кадять вони, але ті помогти не поможуть їм за часу їхнього лиха!
JER|11|13|Бо богів твоїх за числом твоїх міст, Юдо, і за числом вулиць Єрусалиму наставлено жертівників для Молоха, жертівників, щоб кадити Ваалові.
JER|11|14|А ти не молися за цього народа, і благання й молитви за них не здіймай, бо Я не почую за часу того, коли кликати будуть до Мене з-за лиха свого!
JER|11|15|Пощо Моєму коханому в домі Моєму чинити злі заміри? Чи товсті куски і м'ясо посвятне відвернуть від тебе нещастя твоє? Тоді б ти радів!
JER|11|16|Оливка зелена, гарна плодом хорошим, так кликнув Господь твоє ймення. Але з шумом великого вітру огонь запалився круг неї, і галузки її поламаються!
JER|11|17|А Господь Саваот, що тебе посадив, говорив був на тебе лихе за зло дому Ізраїля та дому Юди, що робили собі, щоб гнівити Мене, щоб кадити Ваалові.
JER|11|18|А Господь дав пізнати мені й я пізнав, і тоді Ти вчинив, що побачив я їхні діла.
JER|11|19|А я був, мов лагідна вівця, що провадять її на заколення, і не знав, що на мене вони вимишляли затії: Понищмо це дерево з плодом його, і з краю живих його витнім, і ймення його не згадається більше!
JER|11|20|Але, Господи Саваоте, Ти Суддя справедливий, що досліджуєш нирки та серце, хай над ними побачу я помсту Твою, бо справу свою я довірив Тобі!
JER|11|21|Тому так промовляє Господь на людей Анатоту, що пошукують душу твою та говорять: Не пророкуй Ім'ям Господа, щоб не померти тобі від рук наших!
JER|11|22|Тому так промовляє Господь Саваот: Ось Я навіщу їх: від меча юнаки повмирають, а сини їхні та їхні дочки від голоду вмруть!
JER|11|23|І останку не буде по них, бо спроваджу Я зло на людей Анатоту у році навіщення їх!...
JER|12|1|Справедливий Ти, Господи, будеш, коли б я судився з Тобою, проте правуватися буду з Тобою: чому то дорога безбожним щаститься, чому то спокійні всі зрадники?
JER|12|2|Ти їх посадив і вони вкоренились, ростуть і приносять плоди. Ти близький в устах їхніх, та далекий від їхніх сердець.
JER|12|3|А Ти, Господи, знаєш мене, Ти бачив мене й дослідив моє серце, що з Тобою воно. Відлучи їх, немов на заріз ту отару, і признач їх на день побиття!
JER|12|4|Аж доки в жалобі земля пробуватиме, і сохнути буде трава всього поля за зло її мешканців? Гине худоба та птаство, бо сказали вони: кінця нашого Він не побачить!
JER|12|5|Як ти з пішими бігав, і вони тебе змучили, то як будеш змагатися з кіньми? Ти в спокійному краї безпечний, та що будеш робити в повідді Йордану?
JER|12|6|Бо також твої браття та дім твого батька і вони тебе зраджують, і криком кричать за тобою, не вір їм, коли й добре тобі говоритимуть!
JER|12|7|Покинув Я Свій дім, залишив спадок Свій; миле Моєї душі Я віддав у долоню її ворогів.
JER|12|8|Спадок Мій Мені став, мов лев той у лісі, свій голос дав проти Мене, тому то його Я зненавидив...
JER|12|9|Чи для Мене спадок Мій, хижий птах різнобарвний, що хижі птахи позлітались круг нього? Ідіть, позбирайте усю польову звірину, спровадьте, щоб жерли!
JER|12|10|Численні пастирі попсували Мого виноградника, потоптали Мій уділ, Мій улюблений уділ вони обернули на голу пустиню!
JER|12|11|Обернули його на спустошення, він при Мені у жалобі, спустошений, увесь Край опустілий, бо нікого нема, хто б поклав це на серце собі!
JER|12|12|Поприходять на всі лисі гори в пустині руїнники, бо меч Господа все позжирає від краю землі й аж до краю землі, миру не буде для всякого тіла!...
JER|12|13|Пшеницю посіяли, терня ж пожали, намучилися, та не мали користи... І буде вам сором за ваші плоди через лютість Господнього гніву!
JER|12|14|Так говорить Господь про лихих усіх сусідів моїх, що вони дотикаються того спадку, що Я дав на спадщину народу Моєму Ізраїлеві: Ось Я повириваю їх з їхньої землі, і вирву дім Юдин з середини їхньої.
JER|12|15|І станеться, як Я їх повириваю, то вернуся й помилую їх, і кожного з них приверну до спадщини його, і кожного до краю його.
JER|12|16|І буде, якщо вони справді навчаться доріг народу Мого, щоб присягатися Йменням Моїм: Як живий Господь, як вони присягати навчили народ Мій Ваалом, то збудуються серед народу Мого!
JER|12|17|А якщо не послухають, то вирву народ цей, вириваючи та вигубляючи, каже Господь!
JER|13|1|Так промовив до мене Господь: Іди й купи собі льняного пояса, і підпережи ним свої стегна, але в воду не клади його.
JER|13|2|І купив я того пояса за Господнім словом, та й підперезав свої стегна.
JER|13|3|І було мені слово Господнє удруге, говорячи:
JER|13|4|Візьми того пояса, якого купив, що на стегнах твоїх, і встань, іди до Ефрату, та й сховай його там у розщілині скелі.
JER|13|5|І пішов я, і сховав його в Ефраті, як Господь наказав був мені.
JER|13|6|І сталося по багатьох днях, і сказав мені Господь: Устань, іди до Ефрату, і візьми звідти того пояса, що Я наказав був тобі сховати його там.
JER|13|7|І пішов я до Ефрату, і викопав, і взяв того пояса з місця, де я сховав був його, аж ось той пояс нездатний!
JER|13|8|І було мені слово Господнє, говорячи:
JER|13|9|Так говорить Господь: Отак знищу Я Юдину гордість та гордість велику Єрусалиму,
JER|13|10|цього злого народа, що не хоче він слухатися Моїх слів, що ходить за впертістю серця свого! І пішов він в сліди інших богів, щоб служити їм та поклонятися їм. І станеться він, як цей пояс, до нічого нездатний!...
JER|13|11|Бо як прилягає цей пояс до стегон чоловіка, так притвердив Я до себе ввесь Ізраїлів дім та ввесь Юдин дім, говорить Господь, щоб стали народом Мені і йменням, і хвалою та пишнотою, та вони не послухались!
JER|13|12|І скажеш до них оце слово: Так говорить Господь, Бог Ізраїлів: усякий бурдюк вином наповняється. І відкажуть тобі: Чи ми справді не знаєм, що всякий бурдюк вином наповняється?
JER|13|13|І скажеш до них: Так говорить Господь: Ось наповню Я п'янством усіх мешканців Краю цього, і царів, що сидять на Давидовім троні, і священиків, і пророків, і всіх мешканців Єрусалиму.
JER|13|14|І розіб'ю їх одного об одного, разом батьків та синів, говорить Господь, Не змилуюся, і не змилосерджусь, і не пожалію, щоб їх не понищити!
JER|13|15|Послухайте ви та візьміть до ушей, не вивищуйтеся, бо Господь це сказав!
JER|13|16|Дайте Господу, Богові вашому, славу, поки не зробить Він темно, і поки на темних горах не спіткнуться вам ноги! І будете ви сподіватися світла, а Він зробить це темрявою та вчинить імлою...
JER|13|17|А коли ви цього не послухаєте, буде плакати таємно душа моя з вашої гордости, й око моє проливатиме сльози, і зайдеться сльозою, бо стадо Господнє займуть у полон!...
JER|13|18|Скажіть до царя й до царевої матері: Сідайте додолу, бо з голів ваших спала корона вашої слави!
JER|13|19|Південні міста позамикані будуть, і не буде, хто б їх відчинив, вигнаний буде ввесь Юда, вигнаний буде цілком!
JER|13|20|Зведіть ваші очі, й побачте отих, що приходять із півночі: де череда та, що дана тобі, отара пишноти твоєї?
JER|13|21|Що ти скажеш, о дочко Сіону, як Він над тобою панами поставить отих, яких ти навчила була за довірених бути, чи ж муки не схоплять тебе, немов ту породіллю?
JER|13|22|коли ж скажеш у серці своєму: Чому такі речі спіткали мене? за численні провини твої відкриті подолки твої, оголені ноги твої силоміць!
JER|13|23|Чи мурин відмінить коли свою шкіру, а пантера ті плями свої? Тоді зможете й ви чинити добре, навчені чинити лихе!
JER|13|24|Тому розпорошу їх, мов ту полову, що з вітром з пустині летить:
JER|13|25|Оце жеребок твій, це уділ, який Я відміряв тобі, говорить Господь, бо забула Мене та надіялася на неправду!
JER|13|26|І закочу теж подолки твої над обличчя твоє, і покажеться ганьба твоя:
JER|13|27|твої перелюбства й іржання твої, сором блуду твого на полі на пагірках, Я бачив гидоти твої... Горе тобі, Єрусалиме, що не очистишся! Доки ж іще?
JER|14|1|Слово Господнє до Єремії, що було в справі посухи.
JER|14|2|Упала в жалобу Юдея, а брами її ослабіли, насупилися на землі, і знявся крик Єрусалиму.
JER|14|3|А вельможі її своїх слуг посилають по воду, вони йдуть до криниці й води не знаходять, їхній посуд порожній вертається... Засоромляться та зашаріють вони, і свої голови понакривають.
JER|14|4|Тому, що земля стала спрагла, бо дощу не було на землі, засоромилися рільники, свої голови понакривали.
JER|14|5|Навіть ланя на полі породить сарнятко та й кине, бо немає трави...
JER|14|6|Навіть дикі осли поставали на голих горах, вітер втягують, мов ті шакали, і меркнуть їм очі, бо немає трави...
JER|14|7|Якщо проти нас свідчать наші провини, о Господи, то зроби ради Ймення Свого, бо намножились наші відступники, ми Тобі нагрішили!
JER|14|8|О надіє Ізраїлева, о Спасителю в часі недолі, нащо будеш Ти в Краї, як той чужаниця, й як той подорожній, що намета лише на ночліг розтягає?
JER|14|9|Нащо будеш Ти, мов людина остовпіла, немов той силач, що не може спасти? Таж Ти в нашій середині, Господи, Ймення ж Твоє на нас кличеться, не залишай нас!
JER|14|10|Так говорить Господь до народу цього: Так люблять вони волочитись, а не стримувати своїх ніг, тому то не має Господь уподобання в них, Він тепер їхню провину згадає, і їхній гріх покарає!
JER|14|11|І промовив до мене Господь: Не молись за народ цей на добре йому:
JER|14|12|Як вони будуть постити, Я не послухаю їхніх благань, а коли принесуть цілопалення й дар, Я їх не прийму, бо Я повигублюю всіх їх мечем, і голодом, і моровицею!...
JER|14|13|А я відказав: О Господи, Боже! Ось пророки говорять до них: Ви не будете бачити меча, і не буде вам голоду, правдивий бо мир в цьому місці вам дам!
JER|14|14|Та промовив до мене Господь: Ці пророки неправду Іменням Моїм пророкують: Я їх не посилав, і не наказував їм, і їм не говорив! Вони вам пророкують невірні видіння та чари, нікчемність й оману свого серця...
JER|14|15|Тому так промовляє Господь на пророків, які пророкують Іменням Моїм, хоч Я не посилав їх, та що кажуть вони: Меч та голод не буде в цім Краї: від меча та від голоду згинуть пророки такі!
JER|14|16|А народ, що таке пророкують йому, розкиданий буде по вулицях Єрусалиму від голоду та від меча, і не буде кому поховати його, вони й їхні жінки, й їхні сини та їхні дочки, і виллю на них їхнє зло!
JER|14|17|І ти скажеш до них оце слово: Хай заходять удень та вночі мої очі слізьми, і нехай не затихнуть, бо дівчина, доня народу мого, буде побита великим нещастям, дуже болючим ударом!
JER|14|18|Якщо вийду на поле ось побиті мечем, й якщо вийду до міста ось помлілі із голоду, і навіть пророк та священик шмигляють по краю, якого не знають...
JER|14|19|Чи насправді покинув Ти Юду? Чи й Сіоном гидує душа Твоя? Чому вразив Ти нас і немає нам ліку? Ми чекаємо миру й немає добра, і часу вздоровлення та ось тільки жах!...
JER|14|20|Знаємо, Господи, нашу безбожність, вину наших батьків, бо ми проти Тебе згрішили,
JER|14|21|та не відкидай нас ради Ймення Свого, не безчесть трону слави Своєї, пам'ятай, не зламай заповіту Свого із нами!
JER|14|22|Хіба є між марними божками поганів такі, що спускають дощі? І чи небо саме дає зливу? Чи ж не Ти Господь Бог наш? Тому то на Тебе надіємось ми, бо Ти це все чиниш!
JER|15|1|І промовив до мене Господь: Якщо став би Мойсей й Самуїл перед лицем Моїм, то душа Моя до народу цього не звернулася б! Віджени їх із-перед Мого лиця, і нехай повиходять!
JER|15|2|І буде, як скажуть до тебе вони: Куди підемо? то скажеш до них: Так говорить Господь: Хто на смерть ті на смерть, і хто на меча на меча, і хто на голод на голод, а хто до полону в полон...
JER|15|3|І Я навіщу їх чотирьома способами, говорить Господь: мечем, щоб побити, і псами, щоб їх волочити, і птаством небесним, і земною звіриною, щоб жерли та нищили...
JER|15|4|І Я дам їх на пострах усім царствам землі за Манасію, Єзекіїного сина, царя Юдиного, за те, що зробив був він в Єрусалимі.
JER|15|5|Бо хто змилується над тобою, о Єрусалиме? І хто співчуття тобі виявить? І хто зверне з путі, щоб тебе запитати про поводження?
JER|15|6|Ти покинув Мене, промовляє Господь, відступився назад, тому Я простягнув Свою руку на тебе, і знищив тебе, утомився Я жалувати!
JER|15|7|І віячкою їх розвіяв по брамах землі, позбавив дітей, і погубив Свій народ, бо вони не вернулись з доріг неправдивих своїх,
JER|15|8|у Мене більше було його вдів, як морського піску! А на матір юнацтва, спровадив опівдні грабіжника їм, нагло кинув на неї страхіття та жах,
JER|15|9|зомліла вона, що сімох породила, видихнула свою душу, зайшло сонце її, коли був іще день, засоромилася та збентежилась... А решту їх Я дам під меча перед їхніми ворогами, говорить Господь...
JER|15|10|Горе мені, моя мати, що ти породила такого мене, чоловіка сварливого та чоловіка сутяжного для всієї землі! Нікому я не позичав, і ніхто мені не боргував, та всі проклинають мене...
JER|15|11|Промовив Господь: Я справді підсилю на добре тебе, Я справді вчиню, що проситиме ворог тебе за час зла й за час утиску!
JER|15|12|Чи можна зламати залізом залізо із півночі й мідь?
JER|15|13|Багатство твоє й твої скарби на здобич віддам, і не за ціну, але за гріхи твої всі, у всіх границях твоїх.
JER|15|14|І вчиню, що ти будеш служити своїм ворогам у тім краї, якого не знаєш, бо огонь запалав в Моїм гніві, і над вами палатиме він!
JER|15|15|Ти, Господи, знаєш усе, згадай же мене й заступися за мене, і помстися над тими, що гонять мене! На довгу Свою терпеливість до них мене не бери, знай, що сором носив я за Тебе!
JER|15|16|Як тільки слова Твої знаходилися, то я їх поїдав, і було слово Твоє мені радістю і втіхою серця мого, бо кликалось Ймення Твоє надо мною, о Господи, Боже Саваоте!
JER|15|17|Не сидів я на зборі веселому та не радів, через руку Твою я самітний сидів, бо Ти гнівом наповнив мене.
JER|15|18|Чому біль мій став вічний, а рана моя невигойна, що не хоче загоїтись? Чи справді Ти станеш мені як обманний потік, що води його висихають?
JER|15|19|Тому Господь так відказав: Якщо ти навернешся, то тебе приверну, і перед лицем Моїм станеш, а як здобудеш дорогоцінне з нікчемного, будеш як уста Мої: до тебе самі вони звернуться, а не ти до них звернешся!
JER|15|20|І дам Я тебе для оцього народу за мура міцного із міді, і будуть вони воювати з тобою, та не переможуть тебе: бо Я буду з тобою, щоб спасати тебе й щоб тебе рятувати, говорить Господь!
JER|15|21|І врятую тебе з руки злих, і з рук насильників тих тебе визволю!
JER|16|1|І було слово Господнє до мене, промовляючи:
JER|16|2|Не бери собі жінки, і хай у тебе не буде синів, ні дочок у цьому місці.
JER|16|3|Бо так промовляє Господь про синів і про дочок, що народжені в місці цьому, і про їхніх матерів, що народжують їх, і про їхніх батьків, що їх родять у Краї цьому:
JER|16|4|Від жахливих хворіб повмирають вони, не будуть оплакувані, і не будуть поховані, гноєм стануть вони на поверхні землі... Від меча та від голоду згинуть вони, і стане їхній труп стервом птаству небесному й земній звірині...
JER|16|5|Бо так промовляє Господь: Не заходь у дім смутку, і не ходи голосити, і не співчувай їм, бо від цього народу забрав Я Свій мир, говорить Господь, ласку та милість.
JER|16|6|І повимирають великі й малі в цьому Краї, не будуть поховані, і голосити не будуть за ними, і не будуть робити нарізів, і не будуть робити собі лисини...
JER|16|7|І не будуть ламати їм хліба в жалобі, щоб потішити їх над померлим, і не напоять їх келіхом втіхи над батьком його й його матір'ю...
JER|16|8|І до дому бенкету не входь, щоб сидіти із ними, щоб їсти й щоб пити.
JER|16|9|Бо так промовляє Господь Саваот, Бог Ізраїлів: Ось Я припиню в цьому місці на ваших очах і в днях ваших голос радісний й голос веселий, голос молодого та голос молодої!
JER|16|10|І буде, коли перекажеш народові цьому ці слова, то скажуть тобі: За що Господь говорив проти нас все велике це лихо? І яка вина наша, й який то наш гріх, яким ми прогрішилися Господу, Богові нашому?
JER|16|11|І відкажеш до них: За те, що Мене батьки ваші покинули, каже Господь, і пішли за іншими богами і служили їм та поклонялися їм, а Мене полишили й Закона Мого не виконували!
JER|16|12|А ви робите гірше від ваших батьків, і кожен із вас ось іде за упертістю лютого серця свого, щоб Мені не служити...
JER|16|13|Тому викину вас з цього Краю до краю, якого не знали ні ви, ані ваші батьки. І будете там богам іншим служити удень та вночі, бо не дам Я вам милости.
JER|16|14|Тому наступають ось дні, говорить Господь, і не будуть уже говорити: Як живий Господь, що вивів синів Ізраїлевих із краю єгипетського,
JER|16|15|а тільки: Як живий Господь, що вивів синів Ізраїлевих із північного краю, і зо всіх тих країв, куди був розігнав їх... Та Я їх верну на їхню землю, яку Я був дав батькам їхнім.
JER|16|16|Оце Я пошлю по численних рибалок, говорить Господь, і виловлять їх, немов рибу, а потому пошлю по численних мисливців, і повиловлюють їх з усіх гір, і з усякого взгір'я, і зо скельних розщілин.
JER|16|17|Бо очі Мої на всі їхні дороги: вони не сховалися з-перед Мого лиця, і з-перед ока Мого не закрилася їхня провина.
JER|16|18|І найперше Я їм надолужу подвійно за їхню провину й за гріх їхній, за теє, що трупом обриджень своїх збезчестили Край мій, а їхні гидоти спадок Мій переповнили...
JER|16|19|О Господи, сило моя та твердине моя, і захисте мій в день недолі! Поприходять до тебе народи від кінців землі та й промовлять: Одідичили наші батьки лиш неправду й марноту, пожитку ж від них не було...
JER|16|20|Чи зробить людина для себе богів, а вони не боги?
JER|16|21|Тому то ось Я учиню, що познають цим разом вони, учиню, що познають вони Мою руку та силу Мою, і познають, що Ймення Моє це Господь!
JER|17|1|Гріх Юдин написаний рильцем залізним, діямантовим вістрям він виритий на таблиці їхнього серця, і на рогах жертовників їхніх.
JER|17|2|Як про синів своїх, так пам'ятають про жертовники своїх та своїх Ашер при зеленому дереві, на високих підгірках,
JER|17|3|про гору на полі. Багатство твоє й твої скарби на здобич віддам, пагірки жертовні твої за гріх по всіляких границях твоїх.
JER|17|4|І опустиш ти руку свою спадку свого, що Я дав був тобі... І вчиню, що ти будеш служити своїм ворогам у тім краї, якого не знаєш, бо огонь запалили ви в гніві Моїм, й аж навіки палатиме він!
JER|17|5|Так говорить Господь: Проклятий той муж, що надію кладе на людину, і робить раменом своїм слабу плоть, а від Господа серце його відступає!
JER|17|6|І він буде, як голий той кущ у степу, і не побачить, щоб добре прийшло, і він пробуватиме в краї сухому в пустині, у краї солоному та незамешканому...
JER|17|7|Благословенний той муж, що покладається на Господа, що Господь то надія його!
JER|17|8|І він буде, як дерево те, над водою посаджене, що над потоком пускає коріння своє, і не боїться, як прийде спекота, і його листя зелене, і в році посухи не буде журитись, і не перестане приносити плоду!
JER|17|9|Людське серце найлукавіше над все та невигойне, хто пізнає його?
JER|17|10|Я Господь, що досліджує серце, що випробовує нирки, щоб кожному дати згідно з путтю його, за плодом учинків його.
JER|17|11|Куропатва висиджує яйця, яких не принесла, це той, хто багатство набув, та неправдою: він покине його в половині днів своїх, і стане безумним при своєму кінці...
JER|17|12|Трон слави, високий від віку, це місце нашої святині!
JER|17|13|Надіє Ізраїлева, Господи, посоромлені будуть усі, хто Тебе залишає! Ті, що Мене покидають, на піску будуть списані, бо вони покинули Господа, джерело живої води.
JER|17|14|Уздоров мене, Господи, і буду вздоровлений я, спаси Ти мене, і я буду спасений, бо Ти слава моя!
JER|17|15|Ось вони мені кажуть: Де слово Господнє? Нехай воно прийде!
JER|17|16|А я не відтягавсь бути пастирем в Тебе, не жадав злого дня, Ти це знаєш, що виходило з уст моїх, те перед лицем Твоїм явне було.
JER|17|17|Не будь Ти для мене страхіттям, на день зла Ти моє пристановище!
JER|17|18|Бодай посоромились ті, хто мене переслідує, а я щоб не був посоромлений, нехай побентежені будуть вони, а я хай не буду збентежений, день злого на них наведи та зламай їх подвійним зламанням!
JER|17|19|Так промовив до мене Господь: Іди, і станеш у брамі синів народу, що юдські царі входять нею та нею виходять, та по всіх брамах Єрусалиму.
JER|17|20|І скажеш до них: Послухайте слова Господнього, царі юдські й уся Юдеє, та всі мешканці Єрусалиму, що входите брамами тими.
JER|17|21|Так говорить Господь: Стережіться за душі свої, і не носіть тягару за суботнього дня, і не носіть його брамами Єрусалиму.
JER|17|22|І не носіть тягару з домів ваших суботнього дня, і жодної праці робити не будете, і день суботній освятите, як Я вашим батькам наказав був!
JER|17|23|Та вони не послухали, й вуха свого не схилили, і вчинили себе тугошиїми, щоб не слухатися та не брати навчання.
JER|17|24|І буде, якщо Мене справді ви будете слухатись, каже Господь, щоб тягару не носити в брами міста цього за суботнього дня, і щоб освятити день суботній, і щоб жодної праці в цей день не робити,
JER|17|25|то ходитимуть брамами міста цього царі та князі, що будуть сидіти на троні Давидовім, що їздити будуть колесницями й кіньми, вони й їхні правителі, юдеї та мешканці Єрусалиму, і це місто стоятиме вічно!
JER|17|26|І будуть приходити з Юдиних міст та з околиць Єрусалиму, і з краю Веніяминового, і з рівнини, і з гір, і з півдня, і цілопалення й жертви приносити будуть, та жертву хлібну, і ладан, і будуть приносити жертву подяки до дому Господнього.
JER|17|27|А якщо ви Мене не послухаєтесь, щоб святити день суботній і щоб тягару не носити, і щоб брамами Єрусалиму суботнього дня не ходити, то огонь підпалю в їхніх брамах, і він поїсть єрусалимські палати, і не погасне!
JER|18|1|Оце слово, що було до Єремії від Господа, говорячи:
JER|18|2|Устань, і зійди до дому ганчара, і там почуєш слова Мої.
JER|18|3|І зійшов я до дому ганчара, аж ось він робить працю на кружалі.
JER|18|4|І в руках ганчара попсулась посудина, яку він із глини робив. І він знову зробив з неї іншу посудину, як сподобалося ганчареві зробити.
JER|18|5|І було мені слово Господнє, говорячи:
JER|18|6|Чи не міг би зробити й Я вам, як ганчар цей, о доме Ізраїлів? каже Господь. Ось як глина в руці ганчара, так в руці Моїй, доме Ізраїля, й ви!
JER|18|7|Я часом кажу про народ та про царство, щоб вирвати його, і щоб розбити та вигубити,
JER|18|8|та коли цей народ, що про нього казав Я, повернеться від свого зла, то пожалую Я щодо того зла, яке думав чинити йому.
JER|18|9|А часом кажу про народ та про царство, щоб його збудувати та щоб посадити,
JER|18|10|та як він зробить зле в Моїх очах, щоб не слухатися Мого голосу, то пожалую щодо того добра, про яке говорив, що вчиню Я його.
JER|18|11|А тепер скажи до юдея й до мешканців Єрусалиму, говорячи: Так говорить Господь: Ось готую лихе проти вас, і задумую задум на вас, верніться ж ви кожен з дороги своєї лихої, і поліпшіть дороги свої й свої вчинки!
JER|18|12|Та вони відказали: Пропало! бо ми будем ходити за своїми думками, і кожен робитиме згідно з упертістю серця свого.
JER|18|13|Тому так промовляє Господь: Поспитайте но ви між народами, чи хто чув, як оце? Страшну річ учинила та діва Ізраїлева!
JER|18|14|Хіба сніг Лівану зійде зо скелі на полі? Чи висохнуть води чужі та холодні, текучі?
JER|18|15|Бо про Мене забув Мій народ: вони кадять марноті, а та робить їм так, що вони на дорогах своїх спотикаються, на давніх путях, щоб ходити стежками, по дорозі невбитій,
JER|18|16|щоб свій Край учинити страхіттям, посміховищем вічним... Кожен, хто буде проходити ним, остовпіє та буде хитати головою своєю...
JER|18|17|Мов вітер зо сходу, розвію Я їх перед ворогом; потилицю, а не обличчя Я їм покажу у день їхнього горя!
JER|18|18|І сказали вони: Ходіть, і обміркуємо заміри на Єремію, бо не згинув Закон у священика, і рада в премудрого, а слово в пророка. Ходіть, і удармо його язиком його власним, і не зважаймо на жодні слова його!
JER|18|19|Послухай мене, о мій Господи, і почуй голос моїх супротивників!
JER|18|20|Хіба замість доброго злим надолужено буде? Бо яму копають вони для моєї душі... Згадай же, що перед обличчям Твоїм я стояв, щоб добре про них говорити, щоб гнів Твій від них відвернути!
JER|18|21|Тому їхніх синів віддай голодові, і міццю меча викинь їх з Краю, і бодай жінки їхні дітей погубили та вдовами стали, а їхні чоловіки хай смертю повбивані будуть, юнаки їхні хай будуть побиті мечем на війні!
JER|18|22|Нехай чується крик з їхніх домів, бо орду Ти зненацька спровадиш на них, бо яму копали вони, щоб схопити мене, і для ніг моїх пастки поставили...
JER|18|23|А Ти, Господи, знаєш увесь їхній замір на мене на смерть, не прости їм провин, а гріха їхнього із-перед обличчя Свого не зітри, і хай перед Тобою спіткнуться вони, зроби поміж ними оце під час гніву Свого!
JER|19|1|Господь сказав так: Іди, і купиш баньку в ганчара, і візьми собі з старших народу та з старших священиків.
JER|19|2|І вийдеш до долини Бен-Гіннома, що при вході до Череп'яної брами, і будеш там оголошувати ті слова, що до тебе Я їх говоритиму.
JER|19|3|І скажеш: Послухайте слова Господнього, царі Юди та мешканці Єрусалиму! Так говорить Господь Саваот, Бог Ізраїлів: Ось Я зло наведу на це місце, так що всякому, хто почує про нього, задзвенить в його вухах!
JER|19|4|Це за те, що вони залишили Мене, і вчинили чужим оце місце, і кадили у ньому для інших богів, що не знали їх ані вони, ні батьки їхні, ані юдейські царі, і кров'ю невинних наповнили місце оце,
JER|19|5|і пагірки побудували Ваалові, щоб палити дітей своїх на огні цілопалення для Ваала, чого не велів Я і не говорив, і що на серце Мені не приходило!
JER|19|6|Тому наступають ось дні, говорить Господь, що не буде вже зватися місце це Тофет і Долина Бен-Гіннома, а тільки Долина Убивства.
JER|19|7|І знищу на місці цьому раду Юдину та Єрусалиму, і впадуть від меча перед їхніми ворогами та від руки тих, хто шукає їхньої душі, і дам падло їхнє на стерво для птаства небесного та для земної звірини...
JER|19|8|І вчиню оце місце страхіттям і посміхом, кожен, хто буде проходити ним, остовпіє й засвище, побачивши всі його врази...
JER|19|9|І вчиню, що вони будуть їсти тіло синів своїх й тіло дочок своїх, і тіло один одного їсти вони будуть в облозі та в утискові, яким будуть тиснути їх вороги їхні та ті, хто буде шукати їхню душу...
JER|19|10|І розіб'єш баньку на очах тих людей, що ходять з тобою,
JER|19|11|та й скажеш до них: Так говорить Господь Саваот: Отак розіб'ю Я народ цей та місто оце, як розбивається посуд ганчарський, що не може вже бути направленим, і будуть ховати у Тофеті через брак місця на погреб...
JER|19|12|Так зроблю цьому місцю, говорить Господь, та мешканцям його, щоб зробити це місто, як Тофет...
JER|19|13|І стануть доми Єрусалиму та доми царів Юди, як місце те Тофет, нечисті усі ті доми, що кадили на їхніх дахах усім небесним світилам, та лили жертви литі для інших богів!
JER|19|14|І прийшов Єремія з Тофету, куди посилав його Господь пророкувати, і став у дворі Господнього дому, і сказав до всього народу:
JER|19|15|Так говорить Господь Саваот, Бог Ізраїлів: Ось спроваджу до міста цього та до всіх його міст усе те лихо, що Я говорив був на нього, бо вчинили вони свою шию твердою, щоб не слухатися Моїх слів!
JER|20|1|І почув Пашхур, Іммерів син, священик, що був старшим наглядачем, начальник Господнього дому, Єремію, що пророкував ці слова.
JER|20|2|І Пашхур набив пророка Єремію, і посадив його у в'язницю, що була в горішній брамі Веніяминовій, що в Господньому домі...
JER|20|3|І сталося наступного дня, і вивів Пашхур Єремію з в'язниці, а Єремія промовив до нього: Не Пашхур Господь дав ім'я тобі, а тільки Маґор-Міссавів.
JER|20|4|Бо так промовляє Господь: Ось Я зроблю тебе жахом для тебе самого та для всіх твоїх приятелів, і вони попадають від меча ворогів своїх, а очі твої будуть бачити це. А всього Юду віддам у руку царя вавилонського, і він нажене їх до Вавилону, і позабиває їх мечем.
JER|20|5|І дам увесь скарб цього міста та ввесь його здобуток, і всю коштовність його, та всі скарби юдських царів, усе це дам у руку їхніх ворогів, і вони пограбують їх, і візьмуть їх та й відведуть їх до Вавилону...
JER|20|6|А ти, Пашхуре, та всі мешканці дому твого підете до полону. І прийдеш ти до Вавилону, і помреш там, і будеш похований ти та всі твої приятелі, яким ти неправдиво пророкував.
JER|20|7|Намовляв мене, Господи, і був я намовлений, Ти взяв міцно мене й переміг! Я став цілий день посміховищем, кожен глузує із мене...
JER|20|8|Бо коли тільки я говорю, то кричу, кличу: Ґвалт! та Грабіж! і так сталося слово Господнє мені цілий день за ганьбу й посміховище...
JER|20|9|І я був сказав: Не буду Його споминати, і не буду вже Йменням Його говорити! І стало це в серці моїм, як огонь той палючий, замкнений у костях моїх, і я змучивсь тримати його й більш не можу!
JER|20|10|Бо чув я обмову численних, ось острах навколо: Розкажіть, донесемо на нього! Кожен муж, який в мирі зо мною, чатує мого упадку та каже: Може буде обманений і переможемо його, і помстимося над ним!
JER|20|11|Та зо мною Господь, як потужний силач, тому ті, хто женеться за мною, спіткнуться та не переможуть! Будуть сильно вони посоромлені, бо робили без розуму, вічний сором їм буде, який не забудеться!
JER|20|12|А Господь Саваот випробовує праведного, бачить нирки та серце. Хай над ними побачу я помсту Твою, бо Тобі я відкрив свою справу!
JER|20|13|Співайте пісні Господеві, усі хваліть Господа, бо спасає Він душу убогого від руки лиходіїв!
JER|20|14|Проклятий той день, коли я народився, день, коли породила мене моя мати, хай благословенний не буде!
JER|20|15|Проклятий той муж, який сповістив мого батька, говорячи: Народилось тобі дитя-хлопець, а тим справді потішив його!
JER|20|16|І бодай стався муж той, немов ті міста, що Господь зруйнував й не пожалував їх, і нехай чує крик він уранці, а лемент військовий у часі полудня,
JER|20|17|за те, що в утробі мене не забив, і тоді була б стала мені моя мати за гріб мій, а утроба її вагітною навіки була б!...
JER|20|18|Чого то з утроби я вийшов, щоб бачити клопіт й скорботу, і нащо кінчаються в соромі ці мої дні?...
JER|21|1|Слово, що було до Єремії від Господа, коли цар Седекія послав був до нього Пашхура, сина Малкійїного, та священика Цефанію, сина Маасеїного, говорячи:
JER|21|2|Звернися, за нас до Господа, бо Навуходоносор, цар вавилонський, воює проти нас. Може Господь зробить з нами за всіма Своїми чудами, і той відійде від нас!
JER|21|3|І сказав Єремія до них: Так скажіть до Седекії:
JER|21|4|Так говорить Господь, Бог Ізраїлів: Ось Я назад оберну військові знаряддя, що в вашій руці, що ви воюєте ними поза муром з вавилонським царем та з халдеями, які облягають вас, і позбираю їх до середини цього міста.
JER|21|5|І буду Я воювати з вами рукою витягненою та сильним раменом, і в гніві, і в люті, і в великому пересерді!
JER|21|6|І вражу мешканців цього міста, і чоловіка, і худобу, від великої моровиці повмирають вони!
JER|21|7|А потому говорить Господь Я віддам Седекію, Юдиного царя, і його рабів, і народ, і врятованих у цьому місті від моровиці, від меча та від голоду в руку Навуходоносора, царя вавилонського, та в руку ворогів їхніх, що шукають їхньої душі, і він ударить їх вістрям меча, не змилується над ними й не змилосердиться, і не матиме любови!
JER|21|8|А цьому народові скажеш: Так говорить Господь: Ось Я даю перед вами дорогу життя й дорогу смерти.
JER|21|9|Хто сидітиме в цьому місті, той помре від меча, і від голоду та від моровиці; а той, хто перейде і прийде до халдеїв, що вас облягають, буде жити, і стане йому душа його за здобич.
JER|21|10|Бо Я обернув лице Своє на це місто на зле, а не на добре, говорить Господь, воно буде дане в руку царя вавилонського, а він спалить його огнем!...
JER|21|11|А домові царя Юди скажи так: Послухайте слова Господнього:
JER|21|12|Доме Давидів, отак промовляє Господь: Судіть вранці суд і рятуйте грабованого від руки переслідника, щоб не вийшла, немов той огонь, Моя лють, і вона запалає за зло ваших учинків, і не буде кому погасити!
JER|21|13|Ось Я проти тебе, мешканко долини, о скеле рівнини, говорить Господь, на вас, що говорите: Хто прийде на нас і хто ввійде в помешкання наші?
JER|21|14|Бо Я покараю вас згідно із плодом ваших учинків, говорить Господь, і огонь запалю в його лісі, і він пожере всі довкілля його!
JER|22|1|Так говорить Господь: Зійди в дім Юдиного царя, і будеш казати там оце слово,
JER|22|2|та й промовиш: Послухай Господнього слова, о царю юдейський, що сидиш на Давидовім троні, ти й раби твої та народ твій, що входите в брами оці.
JER|22|3|Так говорить Господь: Чиніть правосуддя та правду, і рятуйте грабованого від руки гнобителя, чужинця ж, сироту та вдову не гнобіть, не грабуйте, і крови невинної не проливайте на місці цьому!
JER|22|4|Бо коли оце слово насправді ви виконаєте, то ходитимуть брамами дому оцього царі, що будуть сидіти на троні Давида, що їздити будуть колесницями й кіньми, він і раб його та народ його.
JER|22|5|А якщо не послухаєтесь оцих слів, то клянуся Собою говорить Господь: руїною станеться дім цей!
JER|22|6|Бо так промовляє Господь про дім царя Юди: Ти для Мене Ґілеад, щит Лівану, та поправді кажу Я, тебе оберну на пустиню, на міста незаселені!
JER|22|7|І приготую на тебе отих, що руйнують людину та зброю її, і вони твої кедри добірні зітнуть і їх повкидають в огонь!
JER|22|8|І люди численні ходитимуть містом оцим і будуть казати один до одного: Защо Господь зробив так цьому місту великому?
JER|22|9|І відкажуть: За те, що вони покинули заповіта Господа, Бога Свого, і вклонялися іншим богам, і служили їм.
JER|22|10|Не плачте за вмерлим, і не жалкуйте за ним, але плакати плачте за тим, хто відходить в полон, бо вже не повернеться, і не побачить землі, де він народився...
JER|22|11|Бо так промовляє Господь до Шаллума, сина Йосіїного, царя Юдиного, що царював замість Йосії, свого батька, що вийшов із місця цього: Він сюди вже не вернеться!
JER|22|12|Бо помре він у місці, куди його полонили, Краю ж цього не побачить уже...
JER|22|13|Горе тому, хто несправедливістю дім свій будує, а верхні кімнати безправ'ям, хто каже своєму ближньому працювати даремно, і платні його йому не дає,
JER|22|14|що говорить: Збудую собі дім великий, і верхні кімнати широкі! І вікна собі повирубує, й криє кедриною, і малює червоною фарбою.
JER|22|15|Чи ти зацарюєш тому, що в кедрах ти мешкаєш? Чи ж твій батько не їв та не пив? І коли правосуддя та правду чинив він, тоді було добре йому,
JER|22|16|він розсуджував справу нужденного й бідного, й тоді добре було! Чи не це Мене знати? говорить Господь.
JER|22|17|Хіба твої очі та серце твоє не обернені тільки на користь свою, та щоб проливати кров невинну, і щоб гніт та насилля чинити?...
JER|22|18|Тому так промовляє Господь про Єгоякима, Йосіїного сина, царя Юдиного: Не будуть за ним голосити: О мій брате! й О сестро! Не будуть за ним голосити: О пане й О величносте його!
JER|22|19|Поховають його, немов того осла, волочачи та викидаючи геть за брами Єрусалиму...
JER|22|20|Зійди на Ливан та й кричи, і в Башані свій голос подай, і кричи з Аваріму, бо понищені всі твої друзі...
JER|22|21|Говорив Я тобі в час гаразду твого, але ти казала: Не слухатиму! Це дорога твоя від юнацтва твого, бо не слухалась ти Мого голосу...
JER|22|22|Усіх твоїх пастирів буря розкидає, а коханці твої підуть до полону, справді, тоді посоромлена та побентежена будеш за все своє зло!...
JER|22|23|О ти, що сидиш на Ливані, що кублишся в кедрах, як ти будеш стогнати, як болі й дрижання на тебе спадуть, мов на ту породіллю!
JER|22|24|Як живий Я, говорить Господь, коли б був Конія, син Єгоякимів, цар Юдин, печаткою-перснем на правій руці Моїй, справді Я й звідти тебе зірву!
JER|22|25|І дам Я тебе в руку тих, хто шукає твоєї душі, і в руку тих, що боїшся ти їх, і в руку Навуходоносора, царя вавилонського, і в руку халдеїв...
JER|22|26|І кину тебе й твою матір, яка породила тебе, до іншого краю, де ви не зродились, і там ви повмираєте!
JER|22|27|А до Краю, куди вони прагнуть душею своєю вернутись, туди не повернуться!
JER|22|28|Чи муж цей, Конія, це глиняний посуд, погорджений та розпорошений? Хіба він посудина та непотрібна? Чом відкинені він та насіння його, та й закинені в землю, якої не знають?
JER|22|29|О Краю, мій Краю, о Краю, послухай Господнього слова:
JER|22|30|Так говорить Господь: Запишіть людину оцю самітною, мужем, якому не буде щаститись у днях його, бо нікому з насіння його не пощаститься сидіти на троні Давидовім та панувати ще в Юді!
JER|23|1|Горе пастирям тим, що розгублюють та розганяють отару Мого пасовиська, говорить Господь!
JER|23|2|Тому так промовляє Господь, Бог Ізраїлів, про пастирів тих, що пасуть Мій народ: Ви отару Мою розпорошили й їх розігнали, та не наглядали за ними. Ось тому покараю Я вас за лихі ваші вчинки, говорить Господь!
JER|23|3|А Я позбираю останок отари Своєї зо всіх тих країв, куди Я їх повиганяв був, і їх поверну на пасовиська їхні, і вони порозплоджуються та розмножаться.
JER|23|4|І над ними поставлю Я пастирів тих, які пастимуть їх, і не будуть боятися вже й не злякаються, і не будуть загублені, каже Господь!
JER|23|5|Ось дні наступають, говорить Господь, і поставлю Давидові праведну Парость, і Цар зацарює, і буде Він мудрий, і правосуддя та правду в Краю запровадить.
JER|23|6|За днів Його Юда спасеться, Ізраїль же буде безпечний. А це Його Ймення, яким Його кликати будуть: Господь праведність наша.
JER|23|7|Тому наступають ось дні, говорить Господь, і не будуть уже говорити: Як живий Господь, що вивів синів Ізраїлевих із краю єгипетського,
JER|23|8|а тільки: Як живий Господь, що вивів і випровадив насіння дому Ізраїлевого з північного краю, і зо всіх тих країв, куди їх був повиганяв! І осядуть вони на своїй землі.
JER|23|9|Про пророків. Розривається серце моє в моїм нутрі, тріпочуть всі кості мої, я став, як п'яний, як той муж, що по ньому вино перейшло, через Господа й ради святих Його слів...
JER|23|10|Бо земля перелюбниками стала повна, бо через прокляття потрапила в жалобу земля, повисихали в степах пасовиська, бо стався лихим їхній біг, їхня сила це кривда...
JER|23|11|Бо й пророк та священик грішать, їхнє зло Я знайшов теж у домі Своїм, говорить Господь.
JER|23|12|Тому буде для них їхня дорога, мов сковзанка в темряві, вони будуть попхнені й впадуть через неї, бо зло Я спроваджу на них року навіщення їх, говорить Господь...
JER|23|13|А в тих самарійських пророків Я бачив безглуздя, вони пророкували Ваалом собі, і вчинили блудячим народ Мій, Ізраїля!
JER|23|14|А в єрусалимських пророків Я бачив гидоту: перелюбство й ходіння в неправді, і руки злочинців зміцнили вони, щоб ніхто з свого зла не вернувся... Всі вони Мені стали, немов той Содом, а мешканці його, як Гомора...
JER|23|15|Тому так промовляє Господь Саваот про пророків оцих: Ось Я їх полином нагодую, і водою отруйною їх напою, бо від єрусалимських пророків безбожність пішла для всієї землі!
JER|23|16|Так говорить Господь Саваот: Не слухайте слів цих пророків, що вам пророкують, вони роблять безглуздими вас, висловлюють привиди серця свого, а не слово з уст Господніх.
JER|23|17|Вони справді говорять до тих, що Мене ображають: Господь говорив: Мир вам буде! А кожному, хто ходить в упертості серця свого, говорять вони: Зло не прийде на вас!
JER|23|18|А хто ж то стояв на таємній Господній нараді, і бачив та чув Його слово? Хто до слова Його прислухався й почув?
JER|23|19|Ось буря Господня, як лютість, виходить, а вихор крутливий на голову несправедливих впаде...
JER|23|20|Гнів Господній не вернеться, поки не зробить, і поки не виконає Він замірів серця Свого; наприкінці днів зрозумієте добре все це!
JER|23|21|Цих пророків Я не посилав, вони побігли самі, Я їм не говорив, та вони пророкують.
JER|23|22|А якби в Моїй раді таємній стояли вони, то вони об'являли б народові Моєму слова Мої, і їх відвертали б від їхньої злої дороги, та від зла їхніх учинків.
JER|23|23|Чи Я Бог тільки зблизька, говорить Господь, а не Бог і здалека?
JER|23|24|Якщо заховається хто у криївках, то Я не побачу Його? говорить Господь. Чи Я неба й землі не наповнюю? каже Господь.
JER|23|25|Я чув, що говорять пророки, що Йменням Моїм пророкують неправду й говорять: Мені снилося, снилось мені!...
JER|23|26|Як довго це буде у серці пророків, які пророкують неправду, та пророкують оману свого серця?
JER|23|27|Вони замишляють зробити, щоб народ Мій забув Моє Ймення, їхніми снами, які один одному розповідають, як через Ваала забули були їхні батьки Моє Ймення.
JER|23|28|Той пророк, що йому снився сон, нехай розповідає про сон, а з яким Моє слово, хай каже про слово правдиве Моє, що соломі до збіжжя? говорить Господь.
JER|23|29|Хіба слово Моє не таке, як огонь, говорить Господь, і як молот, що скелю розлупує?
JER|23|30|Тому то ось Я на пророків, говорить Господь, що слова Мої крадуть один від одного.
JER|23|31|Ось Я на пророків, говорить Господь, що вживають свого язика, але кажуть: Це мова Господня!
JER|23|32|Оце Я на тих, що сни неправдиві звіщають, говорить Господь, вони розповідають про них та впроваджують в блуд Мій народ своєю неправдою й глумом своїм, хоч Я не посилав їх і їм не наказував, і вони помогти не поможуть народові цьому, говорить Господь....
JER|23|33|А коли запитає тебе цей народ, чи пророк, чи священик, говорячи: Яке то Господнє пророцтво? то скажеш до них: Ви тягар, і Я вас поскидаю, говорить Господь.
JER|23|34|А пророка й священика та той народ, який скаже: Господній тягар, то Я мужа того й його дім покараю!
JER|23|35|Отак скажете ви один одному й кожен до брата свого: Що Господь відповів, й що Господь говорив?
JER|23|36|А про Господній тягар не згадуйте більш, бо кожному слово його стане за тягара, і ви перекрутили б слова Бога Живого, Господа Саваота, нашого Бога.
JER|23|37|Так пророкові скажеш: Що Господь тобі відповів, і Що Господь говорив?
JER|23|38|Якщо ж будете ви говорити: Господній тягар, тому так промовляє Господь: За те, що ви кажете слово оце: Господній тягар, хоч Я посилав до вас, кажучи: Не говоріте Господній тягар,
JER|23|39|тому конче Я вас підійму, немов тягара, та й викину вас і те місто, що дав був Я вам та вашим батькам, від Свого лиця...
JER|23|40|І дам Я на вас сором вічний та вічну ганьбу, що не буде забута!...
JER|24|1|Господь показав мені, і ось два коші фіґ стояли перед храмом Господнім, потому, як Навуходоносор, цар вавилонський, вигнав Єхонію, Єгоякимового сина, царя Юдиного, та правителів Юдських, і майстра, і слюсаря з Єрусалиму, та й привів їх до Вавилону.
JER|24|2|Один кіш фіґи дуже добрі, як фіґи першого врожаю, а один кіш фіґи дуже злі, яких не їдять через їхню непридатність.
JER|24|3|І промовив до мене Господь: Що ти бачиш, Єреміє? А я відказав: Фіґи. Фіґи добрі дуже добрі, а злі дуже злі, яких не їдять через їхню непридатність.
JER|24|4|І було мені слово Господнє, говорячи:
JER|24|5|Так говорить Господь, Бог Ізраїлів: Як фіґи ці добрі, так оберну Я на добре вигнанців Юдиних, яких Я послав із цього місця до краю халдейського.
JER|24|6|І зверну Я Своє око на них на добро, і поверну їх до цього Краю, і збудую їх, а не розіб'ю, і засаджу їх, а не вирву.
JER|24|7|І дам Я їм серце пізнати Мене, що Я Господь. І вони Мені будуть народом, а Я буду їм Богом, бо вони навернуться до Мене всім серцем своїм!
JER|24|8|А як фіґи ті злі, яких не їдять через їхню непридатність, то так говорить Господь: За такого Я дам Седекію, царя Юдиного, і його правителів та решту Єрусалиму, що залишилися в цьому Краї та що сидять у краї єгипетському.
JER|24|9|І дам їх за острах, на зло для всіх царств землі, на ганьбу та за притчу, на глум та на прокляття в усіх тих місцях, куди вижену їх.
JER|24|10|І пошлю на них меча, і голод та моровицю, аж поки не вигублені будуть на землі, яку Я був дав їм та їхнім батькам!...
JER|25|1|Слово, що було до Єремії про ввесь народ Юдин за четвертого року Єгоякима, сина Йосіїного, царя Юдиного це перший рік Навуходоносора, царя вавилонського,
JER|25|2|що його сказав пророк Єремія про ввесь Юдин народ та до всіх мешканців Єрусалиму, говорячи:
JER|25|3|Від тринадцятого року Йосії, Амонового сина, царя Юдиного, і аж до цього дня, це вже двадцять і три роки, було слово Господнє до мене. І говорив я до вас, говорячи пильно, та не слухали ви.
JER|25|4|І посилав Господь до вас усіх Своїх рабів пророків, рано та пізно, та не слухали ви, і не нахилили свого уха, щоб послухати.
JER|25|5|А вони говорили: Верніться кожен зо своєї злої дороги та зо зла ваших учинків, і сидіть на тій землі, яку Господь дав вам та вашим батькам відвіку й аж навіки.
JER|25|6|І не ходіть за іншими богами, щоб служити їм та щоб вклонятися їм, і не гнівіть Мене роботою ваших рук, і Я не вчиню вам лихого.
JER|25|7|Та ви не прислухалися до Мене, говорить Господь, щоб не гнівити Мене чином рук своїх, на зло собі.
JER|25|8|Тому так промовляє Господь Саваот: За те, що ви не слухалися слів Моїх,
JER|25|9|ось Я пошлю й позбираю всі північні роди, говорить Господь, пошлю до Навуходоносора, царя вавилонського, Мого раба, і наведу їх на Край цей, і на мешканців його та на всіх цих народів навколо, і вчиню їх закляттям, і оберну їх на страхіття, і на посміховище, і на вічні руїни.
JER|25|10|І Я вигублю в них голос радісний та голос веселий, голос молодого та голос молодої, гуркіт жорен та світло світильника...
JER|25|11|І стане цей край руїною, спустошенням, а ці народи будуть служити вавилонському цареві сімдесят літ!
JER|25|12|І станеться, як сповниться сімдесят літ, покараю Я вавилонського царя та цей люд, говорить Господь, за їхню провину, та халдейський край, й оберну його на вічне спустошення.
JER|25|13|І спроваджу на цей край всі Мої слова, що Я говорив був проти нього, усе, що написане в цій книзі, що пророкував Єремія про всі народи.
JER|25|14|Бо їх поневолять численні народи та великі царі, і Я надолужу їм за їхнім чином та за ділом їхніх рук.
JER|25|15|Бо так промовляє до мене Господь, Бог Ізраїлів: Візьми з Моєї руки келіха вина цього гніву, і напоїш ним усі народи, до яких посилаю тебе.
JER|25|16|І будуть вони пити, і будуть хитатися, стратять розум через меча, що Я посилаю між них...
JER|25|17|І взяв я келіха з Господньої руки, і напоїв усі народи, до яких Господь висилав мене:
JER|25|18|Єрусалим та міста Юди, і царів його та правителів його, щоб віддати їх на руїну, на страхіття, на посміховище та на прокляття, як цього дня,
JER|25|19|фараона, царя єгипетського, і рабів його, і правителів його, та ввесь його народ,
JER|25|20|і всю мішанину народів Єгипту, і всіх царів краю Уц, і всіх царів филистимського краю, і Ашкелон, і Аззу, і Екрон, і решту Ашдоду,
JER|25|21|Едома й Моава та синів Аммона,
JER|25|22|і всіх царів Тиру, і всіх царів Сидону, і всіх царів островів, що на тому боці моря,
JER|25|23|і Дедана, і Тему, і Буза, і всіх, що волосся довкола стрижуть,
JER|25|24|і всіх царів Арабії, і всіх царів мішаних народів, що пробувають у пустині,
JER|25|25|і всіх царів Зімрі, і всіх царів Еламу, і всіх царів Мідії,
JER|25|26|і всіх царів півночі, близьких та далеких один від одного, і всі царства землі, що на земній поверхні, а цар Шешаху буде пити по них.
JER|25|27|І скажеш до них: Так говорить Господь Саваот, Бог Ізраїлів: Пийте й впивайтеся, і виметуйте, і падайте та не вставайте перед мечем, що Я посилаю між вас.
JER|25|28|І буде, коли не захочуть вони взяти келіха з твоєї руки на пиття, то промовиш до них: Так говорить Господь Саваот: Конче будете пити!
JER|25|29|Бо ось у місті, що там було кликане Ймення Моє, зачинаю чинити лихе, а чи ви не покарані будете? Покарані будете, бо Я кличу меча на всіх мешканців Краю, говорить Господь Саваот!
JER|25|30|А ти пророкувати їм будеш усі ці слова, й до них скажеш: Господь загримить з височини, і з мешкання святого Свого Свій голос подасть! Загримить на оселю Свою, кликне Він, мов чавильники ті винограду, відповість усім мешканцям земним!
JER|25|31|Дійде гомін до краю землі, бо в Господа пря із народами, Він буде судити кожне тіло і несправедливих віддасть їхньому мечеві, говорить Господь.
JER|25|32|Так говорить Господь Саваот: Ось лихо виходить від люду до люду, і буря велика пробудиться з кінців землі,
JER|25|33|і будуть побиті від Господа в день той лежати від краю землі й аж до краю землі: не будуть оплакувані, і не будуть позбирані, і не будуть поховані, гноєм стануть вони на поверхні землі!...
JER|25|34|Ридайте, о пастирі, та голосіть, і валяйтесь у попелі, проводирі ви отари, бо виповнились ваші дні для зарізу, і вас розпорошу, і впадете, немов дорога та посудина!...
JER|25|35|І не матимуть пастирі захисту, а проводирі череди утікання...
JER|25|36|І чути крик пастирів, і лемент тих проводирів череди, бо пустошить Господь їхню череду,
JER|25|37|і попустошені мирні пасовиська через палання Господнього гніву...
JER|25|38|Він покинув, як лев свою пущу, бо стався страхіттям їхній Край через меча гнобителя, і через запал гніву Його...
JER|26|1|На початку царювання Єгоякима, сина Йосіїного, царя Юдиного, було оце слово від Господа, кажучи:
JER|26|2|Так говорить Господь: Стань на подвір'ї Господнього дому, і будеш говорити всім Юдиним містам, що приходять на поклін до Господнього дому, усі ті слова, що Я наказав був тобі, щоб до них говорити, не вбав ані слова.
JER|26|3|Може почують вони, і вернуться кожен зо своєї злої дороги, й Я пожалую щодо зла, яке думаю вчинити їм через злі їхні вчинки!
JER|26|4|І скажеш до них: Так говорить Господь: Якщо ви не будете прислухуватися до Мене, щоб ходити за Законом Моїм, якого Я дав вам,
JER|26|5|щоб прислухуватися до слів Моїх рабів пророків, яких Я посилаю до вас рано та пізно, та не слухали ви,
JER|26|6|то вчиню з оцим домом, як з Шіло, а місто це дам на прокляття для всіх народів землі...
JER|26|7|І чули священики, і пророки, і ввесь народ Єремію, що говорив ці слова в Господньому домі.
JER|26|8|І сталося, як Єремія закінчив говорити все, що наказав був Господь сказати до всього народу, то схопили його священики, і пророки, і ввесь народ, говорячи: Ти конче помреш!
JER|26|9|Нащо пророкував ти Господнім Ім'ям, кажучи: Як Шіло, буде дім цей, а місто це буде зруйноване, так що не буде в ньому мешканця? І зібрався ввесь народ проти Єремії в Господньому домі.
JER|26|10|І почули ці слова Юдині князі, і відійшли з царського дому до дому Господнього, і сіли при вході до нової Господньої брами.
JER|26|11|І сказали священики та пророки до князів та до всього народу, говорячи: Присуд смерти цьому чоловікові, бо він пророкував проти цього міста, як ви чули своїми вухами!
JER|26|12|І сказав Єремія до всіх князів і до всього народу, говорячи: Господь послав мене пророкувати проти цього дому, і проти цього міста всі ті слова, що ви чули.
JER|26|13|А тепер поліпшіть ваші дороги та ваші чини, і слухайтеся голосу Господа, вашого Бога, то пожалує Господь щодо зла, яке говорив був на вас.
JER|26|14|А я ось я в вашій руці: робіть мені як добре, і як правдиве в ваших очах!
JER|26|15|Тільки справді пізнаєте ви, якщо ви вб'єте мене, що ви невинну кров спровадите на себе й на це місто та на мешканців його, бо Господь справді послав мене до вас говорити в ваші вуха всі ці слова.
JER|26|16|І сказали князі та ввесь народ до священиків та до пророків: Цей чоловік не підлягає присуду смерти, бо він говорив до нас Ім'ям Господа, нашого Бога!
JER|26|17|І встали люди зо старших Краю, і сказали до всього збору народу, говорячи:
JER|26|18|Міхей з Мораші пророкував за днів Єзекії, царя Юдиного, і сказав до всього юдейського народу, говорячи: Так говорить Господь Саваот: Сіон, як те поле, заораний буде, а Єрусалим за румовища стане, а гора цього храму підгірками лісу...
JER|26|19|Чи справді забив його Єзекія, цар Юдин, та ввесь Юда? Чи ж він не побоявся Господа, і не злагодив Господнього лиця? І Господь пожалував щодо того зла, яке говорив був на них. А ми вчинимо таке велике зло на свої душі?
JER|26|20|І також пророкував був Господнім Ім'ям один чоловік, Урійя, син Шемаї, з Кір'ят-Єаріму, і пророкував проти цього міста та проти цього Краю всі ті слова, як Єремія.
JER|26|21|І почув був слова його цар Єгояким, і всі лицарі його та всі князі; і шукав цар способу забити його. І почув це Урійя, і злякався, й утік прийшов до Єгипту.
JER|26|22|І послав цар Єгояким людей до Єгипту, Елнатана, Ахборового сина, і людей з ним до Єгипту.
JER|26|23|І вони вивели Урійю з Єгипту, і привели його до царя Єгоякима, а той ударив його мечем, а трупа його кинув до гробів простих людей...
JER|26|24|Але рука Ахикама, Шаханового сина, була з Єремією, щоб не дати його в руку народу забити його.
JER|27|1|На початку царювання Єгоякима, сина Йосіїного, царя Юди, було оце слово до Єремії від Господа, кажучи:
JER|27|2|Так сказав був до мене Господь: Зроби собі поворозки та ярма, і надінь їх на шию свою.
JER|27|3|І пошлеш їх до царя Едому, і до царя Моаву, і до царя синів Аммону, і до царя Тиру, і до царя Сидону через послів, що приходять до Єрусалиму до Седекії, царя Юдиного.
JER|27|4|І накажеш їм, щоб до своїх володарів говорили: Так говорить Господь Саваот, Бог Ізраїлів: Так скажете вашим володарям:
JER|27|5|Я вчинив землю й людину, і скотину, що на поверхні землі, Своєю силою великою та витягненим раменом Своїм, і дав її тому, хто сподобався в очах Моїх.
JER|27|6|А тепер Я віддав усі ці землі в руку Навуходоносора, царя вавилонського, раба Мого, а також польову звірину дав Я йому, щоб служила йому.
JER|27|7|І будуть служити всі народи йому та синові його, і синові сина його, аж поки не прийде час також його власному краєві, і поневолять його численні народи та великі царі.
JER|27|8|І станеться, той народ і те царство, що не будуть служити йому, Навуходоносорові, цареві вавилонському, і того, хто не дасть шиї своєї в ярмо вавилонського царя, покараю Я народ цей мечем, і голодом, і заразою, говорить Господь, аж поки не зроблю їм кінця рукою його!
JER|27|9|А ви не прислухайтесь до ваших пророків, і до ваших ворожбитів, і до ваших сновидців, і до ваших знахарів, і до ваших чарівників, що говорять до вас, кажучи: Не служіть вавилонському цареві!
JER|27|10|Бо вони пророкують вам неправду, щоб віддалити вас з вашої землі, і Я вас вижену, і ви погинете.
JER|27|11|А народ, що вкладе свою шию в ярмо вавилонського царя й буде служити йому, то залишу його на його землі, говорить Господь, і він буде її обробляти, і буде сидіти на ній.
JER|27|12|І до Седекії, царя Юдиного, говорив Я згідно з усіма цими словами, кажучи: Вкладіть ваші шиї в ярмо вавилонського царя, і служіть йому та його народові, і будете жити.
JER|27|13|Пощо помрете ти та народ твій від меча, голоду та моровиці, як говорив був Господь про той люд, що не буде служити вавилонському цареві?
JER|27|14|І не прислухуйтеся до слів пророків, що кажуть до вас, говорячи: Не будете служити вавилонському цареві, бо неправду вони вам пророкують.
JER|27|15|Бо Я не посилав їх, говорить Господь, і вони пророкують неправду в Ім'я Моє, щоб Я вигнав вас, і погинете ви та пророки, що вам те пророкують!...
JER|27|16|А до священиків та до всього цього народу говорив я, кажучи: Так говорить Господь: Не прислухуйтеся до слів ваших пророків, що пророкують вам, кажучи: Ось тепер незабаром вертається з Вавилону посуд Господнього дому, бо лжу вони пророкують.
JER|27|17|Не прислухуйтеся до них, служіть цареві вавилонському, то будете жити, нащо буде це місто руїною?
JER|27|18|А якщо вони пророки, і якщо слово Господнє з ними, нехай же просять вони Господа Саваота, щоб не перейшов посуд, позосталий в Господньому домі, і в домі царя Юди, і в Єрусалимі до Вавилону.
JER|27|19|Бо так промовляє Господь Саваот про стовпи, і про море, і про підстави, і про решту посуду, позосталого в цьому місті,
JER|27|20|що не забрав їх Навуходоносор, цар вавилонський, коли виганяв був в неволю Єхонію, Єгоякимового сина, царя Юди, з Єрусалиму до Вавилону, та всіх шляхетних Юди та Єрусалиму.
JER|27|21|Бо так промовляє Господь Саваот, Бог Ізраїлів, про посуд, позосталий в Господньому домі та в домі царя Юди та Єрусалиму:
JER|27|22|До Вавилону буде він спроваджений, і там пробуватиме аж до дня Моїх відвідин їх, говорить Господь, тоді випроваджу його, і верну його до цього місця...
JER|28|1|І сталося того року на початку царювання Седекії, царя Юди, четвертого року, п'ятого місяця, сказав до мене Ананія, син Аззурів, пророк, що з Ґів'ону, у Господньому домі, на очах священиків та всього народу, говорячи:
JER|28|2|Так говорить Господь Саваот, Бог Ізраїлів, кажучи: Зламаю ярмо царя вавилонського!
JER|28|3|За два роки часу Я верну до цього місця ввесь посуд Господнього дому, що забрав був Навуходоносор, цар вавилонський, з цього місця, і спровадив його до Вавилону.
JER|28|4|І Єхонію, Єгоякимового сина, царя Юди, і всіх Юдиних вигнанців, що прийшли до Вавилону, Я верну до цього місця, говорить Господь, бо зламаю ярмо царя вавилонського!
JER|28|5|І говорив пророк Єремія до пророка Ананії на очах священиків і на очах усього народу, що стояли в Господньому домі.
JER|28|6|І сказав пророк Єремія: Амінь! Нехай так зробить Господь, нехай виконає Господь слова твої, що ти пророкував про поворот посуду Господнього дому та всього вигнання в неволю з Вавилону до цього місця.
JER|28|7|Тільки послухай це слово, що я говорю в вуха твої та в вуха всього народу:
JER|28|8|Ті пророки, що від віків були передо мною і перед тобою, пророкували про численні краї та про царства великі, про війни, і про голод та про моровицю.
JER|28|9|Пророк, що пророкує про мир, коли справдиться слово пророче, буде пізнаний цей пророк, що його справді послав Господь.
JER|28|10|І взяв пророк Ананія ярмо з шиї пророка Єремії, і поламав його.
JER|28|11|І сказав Ананія на очах усього народу, говорячи: Так говорить Господь: Отак поламаю ярмо Навуходоносора, царя вавилонського, за два роки часу, з шиї всіх народів! І пішов пророк Єремія своєю дорогою.
JER|28|12|І було слово Господнє до Єремії по тому, як пророк Ананія поламав ярмо з шиї пророка Єремії, говорячи:
JER|28|13|Іди, і скажеш до Ананії, говорячи: Так говорить Господь: Ти поламав дерев'яне ярмо, але Я зроблю замість нього ярмо залізне.
JER|28|14|Бо так промовляє Господь Саваот, Бог Ізраїлів: Я дав на шию всіх цих народів залізне ярмо, щоб вони служили Навуходоносорові, цареві вавилонському, і вони будуть служити йому, і навіть польову звірину віддам Я йому!
JER|28|15|І сказав пророк Єремія до пророка Ананії: Послухай же, Ананіє: Не посилав тебе Господь, але ти доводиш, що народ цей довіряє неправді.
JER|28|16|Тому так промовляє Господь: Ось Я викидаю тебе з поверхні землі, цього року ти помреш, бо про відступство від Господа говорив ти!...
JER|28|17|І помер пророк Ананія того року сьомого місяця...
JER|29|1|А оце слова листа, якого пророк Єремія послав з Єрусалиму до залишку старших, і до священиків, і до пророків, і до всього народу, що його вигнав Навуходоносор з Єрусалиму до Вавилону, в неволю,
JER|29|2|по виході царя Єхонії й матері царя та евнухів, князів Юди та Єрусалиму, і майстрів та слюсарів Єрусалиму,
JER|29|3|через Ел'асу, Шафанового сина, та Ґемарію, сина Хілкійїного, яких послав Седекія, цар Юди, до Навуходоносора, царя вавилонського, до Вавилону, говорячи:
JER|29|4|Так говорить Господь Саваот, Бог Ізраїлів, до всього вигнання в неволю, що Я вигнав з Єрусалиму до Вавилону:
JER|29|5|Будуйте доми, і осядьте, і засадіть садки, і споживайте їхній плід!
JER|29|6|Поберіть жінок, і зродіть синів та дочок, і візьміть для ваших синів жінок, а свої дочки віддайте людям, і нехай вони породять синів та дочок, і помножтеся там, і не малійте!
JER|29|7|І дбайте про спокій міста, куди Я вас вигнав, і моліться за нього до Господа, бо в спокої його буде і ваш спокій.
JER|29|8|Бо так промовляє Господь Саваот, Бог Ізраїлів: Нехай не зводять вас ваші пророки, що серед вас, та ваші чарівники, і не прислухуйтеся до ваших снів, що вам сняться.
JER|29|9|Бо лжу вони вам пророкують Ім'ям Моїм, Я їх не посилав, говорить Господь.
JER|29|10|Бо так промовляє Господь: По сповненні семидесяти літ Вавилону Я до вас завітаю, і справджу Своє добре слово про вас, щоб вернути вас до цього місця.
JER|29|11|Бо Я знаю ті думки, які думаю про вас, говорить Господь, думки спокою, а не на зло, щоб дати вам будучність та надію.
JER|29|12|І ви кликатимете до Мене, і підете, і будете молитися Мені, а Я буду прислуховуватися до вас.
JER|29|13|І будете шукати Мене, і знайдете, коли шукатимете Мене всім своїм серцем.
JER|29|14|І Я дамся вам знайти Себе, говорить Господь, і верну вас, і зберу вас зо всіх народів та зо всіх місць, куди Я вигнав був вас, говорить Господь, верну вас до того місця, звідки вас Я був вигнав.
JER|29|15|Якщо ви кажете: Господь поставив нам пророків і в Вавилоні,
JER|29|16|то так говорить Господь до царя, що сидить на Давидовому троні, та до всього народу, що сидить у цьому місті, до ваших братів, що не вийшли з вами на вигнання:
JER|29|17|Так говорить Господь Саваот: Ось Я пошлю на вас меча, голод та моровицю, і дам їх, як обридливі фіґи, яких не їдять через їхню непридатність.
JER|29|18|І буду гнатися за ними мечем, голодом та моровицею, і дам їх на пострах для всіх земних царств, на прокляття, і на остовпіння, і на посміховище, і на ганьбу серед усіх народів, куди Я їх був повиганяв,
JER|29|19|за те, що не слухалися слів Моїх, говорить Господь, що посилав Я до них рабів Моїх пророків, рано та пізно, та не слухали ви, говорить Господь.
JER|29|20|А ви, все вигнання, що послав Я з Єрусалиму до Вавилону, послухайте слова Господнього:
JER|29|21|Так говорить Господь Саваот, Бог Ізраїлів, про Ахава, сина Колаїного, і про Седекію, сина Маасеїного, що неправду пророкують вам Моїм Ім'ям: Ось Я віддам їх у руку Навуходоносора, царя вавилонського, і він повбиває їх на ваших очах!
JER|29|22|І візьметься від них прокляття для всього Юдиного вигнання, що в Вавилоні, говорячи: Нехай учинить тебе Господь, як Седекію та як Ахава, яких вавилонський цар пік на огні,
JER|29|23|за те, що вони зробили огиду в Ізраїлі, і перелюб чинили з жінками своїх ближніх, і говорили ложне слово Ім'ям Моїм, чого Я не звелів їм, а Я відаю це, і Я свідок цьому, говорить Господь.
JER|29|24|А до Шемаї нехеламітянина скажеш, говорячи:
JER|29|25|Так говорить Господь Саваот, Бог Ізраїлів, кажучи: За те, що ти своїм ім'ям посилав листи до всього народу, що в Єрусалимі, і до священика Цефанії, Маасеїного сина, і до всіх священиків, говорячи:
JER|29|26|Господь тебе дав за священика замість священика Єгояди, щоб бути наглядачем у Господньому домі для кожного чоловіка, що божевільний і що вдає пророка, і даси його до в'язниці, а на шию кайдани надінеш.
JER|29|27|А тепер, чому ти не скартав Єремію з Анатоту, що вдає з себе пророка?
JER|29|28|Бо він послав до нас, до Вавилону, говорячи: Довге воно, вигнання! Будуйте доми, і осядьте, і засадіть садки, і споживайте їхній плід!
JER|29|29|І священик Цефанія прочитав цього листа вголос пророкові Єремії.
JER|29|30|І було слово Господнє до Єремії, говорячи:
JER|29|31|Пошли всьому вигнанню, говорячи: Так говорить Господь про нехеламітянина Шемаю: За те, що вам пророкував Шемая, хоч Я не посилав його, і зробив, щоб ви надіялись на неправду,
JER|29|32|тому так промовляє Господь: Ось Я покараю нехеламітянина Шемаю та насіння його: не буде в нього нікого, хто сидів би серед цього народу, і не побачить він добра, яке Я зроблю для народу Свого, говорить Господь, бо про відступство від Господа говорив він!
JER|30|1|Слово, що було до Єремії від Господа, говорячи:
JER|30|2|Так говорить Господь, Бог Ізраїлів, кажучи: Напиши собі всі ті слова, що тобі говорив Я, до книги.
JER|30|3|Бо приходять ось дні, говорить Господь, і Я верну народ Мій Ізраїлів та Юдин, каже Господь, і верну їх до Краю, що їхнім батькам Я був дав, і вони посядуть його.
JER|30|4|А оце ті слова, що Господь говорив про Ізраїля й Юду:
JER|30|5|Бо так промовляє Господь: Почули ми голос страху, переляку, й немає спокою...
JER|30|6|Запитайте й побачте, чи родить мужчина? Чому ж це Я бачу, що в кожного мужа он руки його на стегнах його, немов у породіллі, і всяке обличчя поблідло?
JER|30|7|Ой горе, бо це день великий, немає такого, як він! А це час недолі для Якова, та з нього він буде врятований!
JER|30|8|І буде в той день, говорить Господь Саваот, поламаю ярмо Я із шиї твоєї, а пута твої розірву, і не будуть чужі поневолювати більше його!
JER|30|9|І будуть служити вони тільки Господеві, Богові своєму, і цареві своєму Давидові, якого поставлю Я їм.
JER|30|10|А ти не лякайся, рабе Мій Якові, каже Господь, і не страшися, Ізраїлю, бо Я ось врятую тебе із далекого краю, і нащадків твоїх з краю їхнього полону! І вернеться Яків, і буде спокійний, і буде безпечний, і не буде того, хто б його настрашив,
JER|30|11|бо Я із тобою, говорить Господь, щоб спасати тебе! Бо зроблю Я кінець всім народам, між якими тебе розпорошив, та з тобою кінця не зроблю, і тебе покараю за правом, бо не полишу тебе непокараним!
JER|30|12|Бо так промовляє Господь: Невилічальна пораза твоя, рана твоя невигойна!
JER|30|13|Немає того, хто б справу твою розсудив для твоєї болячки, нема в тебе ліків таких, щоб над раною м'ясо зросло!
JER|30|14|Забули про тебе всі друзі твої, до тебе вони не звертаються, бо ворожим ударом Я вразив тебе, жорстокою карою за численні провини твої, за те, що зміцніли гріхи твої...
JER|30|15|Чого ти кричиш про поразу свою, про свій біль невигойний? За численні твої беззаконства, за те, що зміцніли гріхи твої, Я зробив тобі це...
JER|30|16|Тому всі, що тебе поїдають, поїджені будуть, а всі вороги твої всі вони підуть в полон, і стануть здобиччю ті, хто тебе обдирає, а всіх, хто грабує тебе, на грабунок віддам!
JER|30|17|Бо вирощу шкурку на рані тобі, і з пораз тебе вилікую, говорить Господь, бо відкинута звано тебе, ти, Сіонська дочка, якої ніхто не шукає.
JER|30|18|Так говорить Господь: Ось Я поверну з полону шатра Яковові, і змилуюся над місцями його пробування, і на пагірку своїм побудується місто, а палац осядеться на відповідному місці своїм.
JER|30|19|І вийде подяка із них та голос радіючих, і Я їх помножу, і не буде їх мало, і прославлю Я їх і не будуть принижені!
JER|30|20|І сини його стануть, як перше, а збір його буде міцний перед лицем Моїм, і Я покараю всіх тих, хто його переслідує!
JER|30|21|І буде із нього Потужний його, і постане Володар його з-поміж нього, й Я наближу Його, й Він підійде до Мене! Бо хто є такий, що наразить життя своє на небезпеку, щоб до Мене наблизитись? каже Господь.
JER|30|22|І станете ви народом Мені, а Я буду вам Богом!
JER|30|23|Ось буря Господня, лютість виходить, а вихор крутливий на голову безбожних упаде.
JER|30|24|Не спиниться полум'я гніву Господнього, поки Свого не зробить, і поки не виконає замірів серця Свого, ви наприкінці днів зрозумієте це!
JER|31|1|Того часу, говорить Господь, для всіх родів Ізраїля стану Я Богом, вони ж Мені стануть народом!
JER|31|2|Так говорить Господь: Знайшов милість в пустині народ, від меча врятований, Ізраїль іде на свій спочин.
JER|31|3|Здалека Господь з'явився мені та й промовив: Я вічним коханням тебе покохав, тому милість тобі виявляю!
JER|31|4|Ще буду тебе будувати й збудована будеш, о діво Ізраїлева! Ти знов приоздобишся в бубни свої, та й підеш у танок тих, хто бавиться,
JER|31|5|на горах самарійських ще будеш садити виноградники, виноградарі будуть садити й споживати законно собі!
JER|31|6|Настане бо день, коли кликати буде сторожа на Єфремових горах: Уставайте, та підемо ми на Сіон, до Господа, нашого Бога!
JER|31|7|Бо так промовляє Господь: Співайте для Якова з радістю, та головою народів утішайтесь! Розголосіть, вихваляйте й скажіть: Спаси, Господи, народ Свій, останок Ізраїлів!
JER|31|8|Ось Я їх приведу із північного краю, і зберу їх із кінців землі, з ними разом сліпий та кульгавий, важка й породілля, сюди повертаються збори великі!
JER|31|9|Вони прийдуть з плачем, та Я їх попроваджу в утіхах. Я їх до потоків води попроваджу прямою дорогою, не спіткнуться на ній, бо Ізраїлеві Я став Отцем, а Єфрем, перворідний він Мій!
JER|31|10|Народи, послухайте слова Господнього, і далеко звістіть аж на островах та скажіть: Хто розсіяв Ізраїля, Той позбирає його, і стерегтиме його, як пастир отару свою!
JER|31|11|Бо Господь викупив Якова, і визволив його від руки сильнішого від нього.
JER|31|12|І вони поприходять, і будуть співати на вершині Сіону, і до добра до Господнього будуть горнутись, до збіжжя, і до виноградного соку, і до оливи, і до молодої дрібної худоби та до товару великого! І стане душа їхня, немов той напоєний сад, і не відчують уже більше стомлення!
JER|31|13|Тоді дівчина тішитись буде в танку, і разом юнацтво та старші, бо Я оберну їхню жалобу на радість, і Я їх потішу, і їх звеселю в їхнім смутку!
JER|31|14|І душу священиків ситістю Я напою, а народ Мій добром Моїм буде насичений, каже Господь!
JER|31|15|Так говорить Господь: Чути голос у Рамі, плач та ридання гірке: Рахиль плаче за дітьми своїми, не хоче потішена бути за діти свої, бо нема їх...
JER|31|16|Так говорить Господь: Стримай голос свій від голосіння, і від сльози свої очі, бо є нагорода для чину твого, говорить Господь, і вони вернуться з краю ворожого!
JER|31|17|І для твого майбутнього є сподівання, говорить Господь, і до границь твоїх вернуться діти твої!
JER|31|18|Добре Я чую Єфрема, як він головою похитує, плачучи: Покарав Ти мене і покараний я, мов теля те ненавчене! Наверни Ти мене і вернуся, бо Ти Господь Бог мій!
JER|31|19|Бо як я навернувся, то каявся, коли ж я пізнав, то вдарив по стегнах своїх... Засоромився я та збентежений був, бо я ганьбу ношу молодощів своїх.
JER|31|20|Чи Єфрем не Мій син дорогий, чи не люба дитина Моя? То скільки Я не говорю проти нього, завжди сильно його пам'ятаю! Тому то за нього хвилюється нутро Моє, змилосерджуся справді над ним, говорить Господь!
JER|31|21|Постав собі дороговкази, стовпи собі порозставляй, зверни своє серце на биту дорогу, якою ти йшла, і вернися, о діво Ізраїлева, вернися до цих своїх міст!
JER|31|22|Аж доки тинятися будеш, о дочко невірна? Господь бо новину створив на землі: жінка спасатиме мужа!
JER|31|23|Так говорить Господь Саваот, Бог Ізраїлів: Оце слово прокажуть іще в краї Юдиному й по містах його, коли Я верну їх: Хай Господь благословить тебе, оселе ти правди, о горо свята!
JER|31|24|І осядуть на ній Юда та міста його разом усі, селяни та ті, хто ходить з отарою.
JER|31|25|Бо напоюю Я душу змучену, і кожну душу скорботну насичую.
JER|31|26|На це я збудився й побачив, і був мені сон мій приємний.
JER|31|27|Ось дні настають, говорить Господь, і засію Ізраїлів дім та дім Юдин насінням людини й насінням скотини.
JER|31|28|І буде, як Я пильнував був над ними, щоб їх виривати та бурити, і щоб руйнувати, і губити, і чинити лихе, так Я попильную над ними, щоб їх будувати й садити, говорить Господь!
JER|31|29|Тими днями не скажуть уже: Батьки їли неспіле, а оскома в синів на зубах!
JER|31|30|бо кожен за власну провину помре, і кожній людині, що їсть недоспіле, оскома впаде їй на зуби!
JER|31|31|Ось дні наступають, говорить Господь, і складу Я із домом Ізраїлевим і з Юдиним домом Новий Заповіт.
JER|31|32|Не такий заповіт, що його з їхніми батьками Я склав був у той день, коли міцно за руку їх узяв, щоб їх вивести з краю єгипетського. Та вони поламали Мого заповіта, і Я їх відкинув, говорить Господь!
JER|31|33|Бо це ось отой Заповіт, що його по цих днях складу з домом Ізраїля, каже Господь: Дам Закона Свого в середину їхню, і на їхньому серці його напишу, і Я стану їм Богом, вони ж Мені будуть народом!
JER|31|34|І більше не будуть навчати вони один одного, і брат свого брата, говорячи: Пізнайте Господа! Бо всі будуть знати Мене, від малого їхнього й аж до великого їхнього, каже Господь, бо їхню провину прощу, і не буду вже згадувати їм гріха!
JER|31|35|Так говорить Господь, що сонце дає вдень на світло, і порядок місяцеві й зорям на світло вночі, що порушує море й шумлять його хвилі, Господь Саваот Йому Ймення!
JER|31|36|Як відійдуть устави ці з-перед обличчя Мого, говорить Господь, то й насіння Ізраїлеве перестане народом бути перед обличчям Моїм по всі дні.
JER|31|37|Так говорить Господь: Так як небо вгорі незміриме, і не будуть досліджені долі основи землі, то так не відкину і Я все насіння Ізраїлеве за все те, що зробили, говорить Господь!
JER|31|38|Ось дні настають, говорить Господь, і збудується місто оце Господеві від башти Хананеїла аж до брами Наріжної.
JER|31|39|І піде мірничий шнурок той ще далі, прямо аж до Ґареву, й обернеться він до Ґої.
JER|31|40|І долина вся трупів та попелу, і всі поля аж до долини Кедрону, аж до рогу Кінської брами на схід, усе це буде святість для Господа, не знищиться та не зруйнується ввіки вона!
JER|32|1|Слово, що було до Єремії від Господа за десятого року Седекії, царя Юдиного, це вісімнадцятий рік Навуходоносора.
JER|32|2|А тоді військо вавилонського царя облягало Єрусалим, а пророк Єремія був ув'язнений в подвір'ї в'язниці, що була при домі царя Юдиного,
JER|32|3|що ув'язнив його Седекія, цар Юдин, говорячи: Нащо ти пророкуєш отак: Так говорить Господь: Ось Я видам це місто в руку вавилонського царя, і він здобуде його...
JER|32|4|А Седекія, цар Юдин, не втече від руки халдеїв, бо конче буде він даний в руку вавилонського царя, і будуть говорити уста його з його устами, а очі його будуть бачити очі його...
JER|32|5|І заведе він Седекію до Вавилону, і він буде там, аж поки Я відвідаю його, говорить Господь. Коли ж будете воювати з халдеями, не пощаститься вам...
JER|32|6|А Єремія відказав: Було мені слово Господнє таке:
JER|32|7|Ось Ганамеїл, син Шаллума, твого дядька, іде до тебе сказати: Купи собі моє поле, що в Анатоті, бо ти маєш викупне право купити.
JER|32|8|І прийшов до мене Ганамеїл, син дядька мого, за Господнім словом, до подвір'я в'язниці, та й сказав мені: Купи моє поле, що в Анатоті, що в Веніяминовому краї, бо твоє право спадщини й твій викуп, купи собі! І пізнав я, що це слово Господнє.
JER|32|9|І купив я це поле від Ганамеїла, сина дядька мого, що в Анатоті, і відважив йому десять і сім шеклів срібла.
JER|32|10|А написав я купчу, і запечатав, і засвідчив свідками, та й зважив срібло вагою.
JER|32|11|І взяв я купчого листа запечатаного, за законом та уставами, і відкритого.
JER|32|12|І дав я купчого листа Барухові, синові Нерійї, Махсеїного сина, на очах сина дядька мого Ганамеїла та на очах свідків, що написані в купчому листі, на очах усіх юдеїв, що сиділи в подвір'ї в'язниці.
JER|32|13|І наказав я Барухові на їхніх очах, говорячи:
JER|32|14|Так говорить Господь Саваот, Бог Ізраїлів: Візьми ці листи, цього купчого листа, і запечатаного, і того листа відкритого, і даси його в глиняний посуд, щоб заховались на довгий час.
JER|32|15|Бо так промовляє Господь Саваот, Бог Ізраїлів: Ще будуть купуватися доми та поля й виноградники в цьому Краї!
JER|32|16|І молився я до Господа потому, як дав був купчого листа Барухові, Нерейїному синові, промовляючи:
JER|32|17|О Господи, Боже! Ти небо та землю створив Своєю потужною силою та Своїм витягненим раменом, нічого для Тебе нема неможливого!
JER|32|18|Милість Ти тисячам чиниш, і за провину батьків після них віддаєш в лоно їхніх синів, Боже великий та могутній, Господь Саваот Йому Ймення!
JER|32|19|Великий в пораді й могутній у чинах, що очі Твої відкриті на всі дороги людських синів, щоб кожному дати згідно з його дорогою та згідно з плодом його чинів,
JER|32|20|що знаки та чуда чинив Ти в єгипетськім краї, і чиниш їх аж по цей день, і між Ізраїлем, і між народом, і зробив Собі Ймення, як цього дня!
JER|32|21|І Ти вивів народ Свій Ізраїля з краю єгипетського знаками та чудами, і рукою потужною, і раменом витягненим та страхом великим.
JER|32|22|І дав Ти їм Край цей, який їхнім батькам заприсяг був, щоб дати їм Край цей, що тече молоком він та медом.
JER|32|23|І прийшли, і посіли його, та не слухалися Твого голосу, і Законом Твоїм не ходили; усього, що Ти наказав їм робити, вони не робили, і Ти вчинив, що спіткало їх все оце лихо...
JER|32|24|Ось доходять до міста вали, щоб здобути його, й місто віддане буде у руку халдеїв, що воюють із ним, через меч, і голод, і моровицю... І що говорив Ти, стається, і ось Ти це бачиш.
JER|32|25|А Ти ж був сказав мені, Господи Боже: Купи собі поле за срібло, і засвідч купівлю свідками. ось місто віддане буде у руку халдеїв...
JER|32|26|І було Господнє слово до Єремії, говорячи:
JER|32|27|Ось Я Господь, Бог кожного тіла: чи для Мене є щось неможливе?
JER|32|28|Тому так промовляє Господь: Ось Я віддам оце місто у руку халдеїв і в руку Навуходоносора, царя вавилонського, і він здобуде його!
JER|32|29|І прийдуть халдеї, що воюють з цим містом, і підпалять це місто огнем, та й спалять його й ті доми, що приносились жертви Ваалові на їхніх дахах, і лилися литі жертви для інших богів, щоб Мене прогнівити...
JER|32|30|Бо сини Ізраїлеві та сини Юдині тільки зло учиняли на очах Моїх від юнацтва свого, сини бо Ізраїлеві лиш гнівили Мене чином рук своїх, каже Господь...
JER|32|31|Бо місто це стало Мені на Мій гнів та на лютість Мою з того дня, як його збудували, та аж до дня цього, щоб відкинути його від Мого лиця
JER|32|32|за все те зло синів Ізраїлевих та синів Юдиних, яке учинили, щоб гнівити Мене, вони, їхні царі, князі, їхні священики й їхні пророки, і юдеяни й мешканці Єрусалиму...
JER|32|33|І вони обернулись до Мене потилицею, а не обличчям, хоч Я їх навчав рано й пізно, та не слухалися, щоб прийняти науку...
JER|32|34|І поклали гидоти свої в тому храмі, в якому Ім'я Моє кликалося, щоб його занечистити...
JER|32|35|І побудували жертовні пагірки Ваалові, що в долині Бен-Гіннома, щоб через огонь переводити синів своїх та своїх дочок Молохові, чого їм не наказував Я, й що не входило в серце Мені, щоб чинити ту гидоту, щоб уводити Юду у гріх.
JER|32|36|Тому так промовляє Господь, Бог Ізраїлів, до міста цього, про яке ви говорите: Воно віддане буде у руку царя вавилонського мечем, і голодом, і моровицею:
JER|32|37|Ось Я їх позбираю зо всіх тих країв, куди вигнав був їх Своїм гнівом та люттю Своєю й великим Своїм пересердям, і верну їх до місця цього, і посаджу їх безпечно,
JER|32|38|і вони Мені стануть народом, а Я буду їм Богом!
JER|32|39|І дам Я їм серце одне та дорогу одну, щоб боялись Мене по всі дні на добро собі й синам їхнім по них.
JER|32|40|І складу з ними вічного заповіта, що не відвернуся від них, щоб їм не чинити Свого добра, і дам їм у серце Свій страх, щоб не відступали від Мене!
JER|32|41|І буду Я тішитись ними, щоб чинити їм добро, і їх посаджу на землі цій у правді усім Своїм серцем та всією душею Своєю.
JER|32|42|Бо так промовляє Господь: Як спровадив був Я все велике це зло на народ цей, так спроваджу на них все добро, яке провіщав Я про них!
JER|32|43|І купуватимуть поле в цім Краї, про якого ви кажете: Він спустошення, так що немає людини й скотини, він відданий в руку халдеїв.
JER|32|44|І будуть вони купувати поля за срібло, і писати про це у листі, й запечатувати, і свідчити свідками, у краї Веніяминовому та в околицях Єрусалиму, і в містах Юдиних, і в містах гірських, і в містах долішніх, і в містах південних, бо верну їх із полону, говорить Господь!
JER|33|1|І було Єремії Господнє слово вдруге, коли він ще замкнений був на подвір'ї в'язниці, говорячи:
JER|33|2|Так говорить Господь, що чинить оце, Господь, що вформовує це, щоб поставити міцно оце, Господь Його Ймення:
JER|33|3|Покликуй до Мене і тобі відповім, і тобі розповім про велике та незрозуміле, чого ти не знаєш!
JER|33|4|Бо так промовляє Господь, Бог Ізраїлів, про доми цього міста й про доми царів Юди, що їх поруйновано на оборонні вали,
JER|33|5|приходять вони воювати з халдеями, щоб доми понаповнювати людськими трупами, що вразив Я гнівом Своїм та люттю Своєю, і сховав Я від міста оцього обличчя Своє за все їхнє зло:
JER|33|6|Ось Я йому вирощу шкурку на рані, й дам ліки, та їх уздоровлю, і відкрию багатство спокою та правди для них!
JER|33|7|І Я поверну долю Юди, і долю Ізраїля, і їх розбудую, немов напочатку.
JER|33|8|І очищу Я їх з їхньої провини всілякої, що нагрішили Мені, і пробачу всі їхні провини, якими нагрішили Мені, та відпали від Мене.
JER|33|9|І Єрусалим Мені стане за радісне ймення, за хвалу та пишноту всім людям землі, що почують про все те добро, що зробив Я для них! І вони полякаються та затремтять через все те добро та ввесь спокій, який Я для нього вчинив!
JER|33|10|Так говорить Господь: Ще буде почутий на місці оцьому, про яке ви говорите: Воно поруйноване, так що немає людини й немає скотини, у містах Юди й на вулицях Єрусалиму, спустошених так, що немає людини, й немає мешканця, й немає скотини,
JER|33|11|радісний голос та голос веселий, голос молодого та голос молодої, голос тих, що говорять: Хваліть Господа Саваота, бо добрий Господь, бо навіки Його милосердя! що жертву хвали до Господнього дому приносять, бо Я поверну долю Краю цього, як було напочатку, говорить Господь!
JER|33|12|Так говорить Господь Саваот: Ще буде на місці оцьому спустошеному, що немає нічого воно від людини та аж до скотини, та по містах його всіх ще буде пасовисько для пастухів, куди приведуть вони череду на відпочинок!
JER|33|13|У містах у горішніх, у містах долішніх, і в південних містах, і в Веніяминовому краї, і в околицях Єрусалиму, і в містах Юдиних ще проходитиме череда через руки рахуючого, говорить Господь!
JER|33|14|Ось дні настають, говорить Господь, і Я виповню добре те слово, що Я провіщав про Ізраїлів дім і про дім Юдин:
JER|33|15|тими днями та часу того Я Давидові зрощу Пагінця справедливости, Він буде чинити на землі правосуддя та правду!
JER|33|16|Юда буде спасений в тих днях, а Єрусалим буде жити безпечно, і його будуть кликати так: Господь наша правда!
JER|33|17|Бо так промовляє Господь: Нема переводу Давидовим мужам, що мають сидіти на троні дому Ізраїлевого,
JER|33|18|і нема переводу в Левитів священиків перед обличчям Моїм тому мужеві, що буде приносити цілопалення, і спалювати хлібну жертву, і приносити жертву всі дні!
JER|33|19|І було слово Господа до Єремії таке:
JER|33|20|Так говорить Господь: Якщо знищите ви заповіта Мого щодо дня та Мого заповіта щодо ночі, щоб не було дня та ночі в їхньому часі,
JER|33|21|то знищений буде також заповіт Мій з Давидом, рабом Моїм, щоб він сина не мав, який не царював би на троні його, і з Левитами-священиками, слугами Моїми!
JER|33|22|І як незчисленні ті зорі небесні, а морський пісок незміренний, так помножу насіння Давида, Мого раба, та Левитів, що служать Мені!
JER|33|23|І було слово Господа до Єремії таке:
JER|33|24|Хіба ж ти не завважив, як народ цей казав був, говорячи: Обидва ті роди, яких Господь вибрав, відкинув Він їх? І народом Моїм вони нехтують, наче б не був він уже перед ними народом.
JER|33|25|Так говорить Господь: Якщо заповіта Мого щодо дня та щодо ночі нема, якщо Я уставів для неба й землі не поклав,
JER|33|26|то відкину й насіння Якова та раба Мого Давида, щоб не брати володарів із насіння його для насіння Авраама, Ісака та Якова... Та не буде того, бо верну їхню долю, й помилую їх!
JER|34|1|Слово, що було Єремії від Господа, коли Навуходоносор, цар вавилонський, і все військо його, і всі царства землі, панування руки його, та всі народи воювали проти Єрусалиму та проти всіх міст його, кажучи:
JER|34|2|Так говорить Господь, Бог Ізраїлів: Іди, і скажеш до Седекії, царя Юдиного, і звістиш йому: Так говорить Господь: Ось Я віддам оце місто в руку вавилонського царя, та й спалю його огнем.
JER|34|3|А ти не втечеш із руки його, бо справді будеш схоплений ти, і в руку його будеш відданий, і очі твої побачать очі вавилонського царя, і уста його говоритимуть з устами твоїми, і до Вавилону ти прийдеш.
JER|34|4|Але послухай Господнього слова, Седекіє, царю Юдин: Так про тебе говорить Господь: Не помреш від меча!
JER|34|5|У мирі помреш ти; і як палили на погребі батькам твоїм, першим царям, що були перед тобою, так будуть палити й тобі, й О пане будуть голосити тобі, бо Я говорив тобі слово, каже Господь.
JER|34|6|І говорив пророк Єремія до Седекії, царя Юдиного, всі оці слова в Єрусалимі.
JER|34|7|А військо вавилонського царя воювало з Єрусалимом та зо всіма позосталими містами Юдиними, з Лахішем та з Азекою, бо вони залишилися серед Юдиних міст містами твердинними.
JER|34|8|Слово, що було до Єремії від Господа по тому, як цар Седекія склав був заповіта з усім народом, що в Єрусалимі, щоб оголосити їм волю,
JER|34|9|щоб кожен відпустив раба свого, і кожен свою невільницю, єврея та єврейку, вільними, щоб ніхто не поневолював свого брата юдея.
JER|34|10|І послухалися всі князі та ввесь народ, що пристали до заповіту, щоб кожен відпустив свого раба, і кожен свою невільницю, вільними, щоб більш не неволити їх. І вони послухалися, і повідпускали.
JER|34|11|Але потому вони знову вернули тих рабів та тих невільниць, яких повідпускали були вільними, і примусили їх стати за рабів та невільниць.
JER|34|12|І було слово Господнє до Єремії від Господа, кажучи:
JER|34|13|Так говорить Господь, Бог Ізраїлів: Я склав був заповіта з вашими батьками того дня, коли виводив їх із єгипетського краю, з дому рабства, кажучи:
JER|34|14|З кінцем семи років відпустите кожен свого брата єврея, що буде проданий тобі й послужить тобі шість років, і відпустиш його вільним від себе. Та не слухалися Мене ваші батьки, і не прихилили свого уха до цього.
JER|34|15|А сьогодні вернулися ви та й зробили справедливе в очах Моїх, щоб оголосити волю кожен своєму ближньому, і склали заповіта перед лицем Моїм у тому домі, в якому кликалось Ім'я Моє.
JER|34|16|Та ви знову збезчестили Ім'я Моє, і вернули кожен раба свого й кожен невільницю свою, яких відпустили були на волю, і примусили їх, щоб були вам рабами та невільницями.
JER|34|17|Тому так промовляє Господь: Ви не послухалися Мене, щоб оголосити волю кожен для брата свого та кожен для свого ближнього, тому то ось Я говорить Господь оголошу вам волю до меча, до моровиці й до голоду, і віддам вас на пострах для всіх царств землі!...
JER|34|18|І віддам цих людей, що переступають Мого заповіта, що не додержують слів заповіту, якого були склали перед лицем Моїм, що вони розрізали надвоє теля та перейшли між його кавалками,
JER|34|19|також князів Юди та князів Єрусалиму, евнухів і священиків, та ввесь народ Краю, що проходили поміж кавалками цього теляти,
JER|34|20|то Я їх віддам у руку їхніх ворогів та в руку тих, хто шукає їхню душу, і стане падло їхнє стервом для птаства небесного та для земної звірини...
JER|34|21|А Седекію, царя Юдиного, та його князів віддам у руку його ворогів та в руку тих, хто шукає їхню душу, та в руку війська вавилонського царя, що відходить від вас.
JER|34|22|Ось Я накажу, говорить Господь, і верну їх до цього міста, і вони воюватимуть з ним, і здобудуть його та й спалять його огнем, а Юдині міста віддам на спустошення, і не буде в них мешканця!...
JER|35|1|Слово, що було до Єремії від Господа за днів Єгоякима, сина Йосії, царя Юди, говорячи:
JER|35|2|Іди до дому Рехавітів, і будеш говорити з ними, і введеш їх до Господнього дому, до однієї з кімнат, і напоїш їх вином.
JER|35|3|І взяв я Яазанію, Єреміїного сина, сина Хаваццініїного, і братів його, і всіх синів його та ввесь дім Рехавітів.
JER|35|4|І ввів я їх до Господнього дому, до кімнати синів Ханана, сина Їґдаліїного, Божого чоловіка, що була при кімнаті князів, що над кімнатою Маасеї, Шаллумового сина, який пильнував порога.
JER|35|5|І поставив я перед синами дому Рехавітів келіхи, повні вина, та чаші, та й сказав до них: Пийте вино!
JER|35|6|А вони відказали: Не будемо пити вина, бо наш батько Йонадав, син Рехавів, наказав нам, говорячи: Не пийте вина ані ви, ані ваші сини аж навіки!
JER|35|7|І не будуйте дому, і не сійте, і не засаджуйте виноградника, і не майте їх, але сидіть у наметах по всі ваші дні, щоб жити довгі дні на поверхні землі, де ви мандруєте!
JER|35|8|І послухалися ми голосу нашого батька Єгонадава, Рехавового сина, про все, що він наказав був нам, щоб не пили вина по всі наші дні ми, наші жінки, наші сини та дочки наші,
JER|35|9|і щоб ні будувати домів для нашого пробування, а виноградник і поле та насіння не будуть наші.
JER|35|10|І осіли ми в наметах, і послухалися, та й зробили все, що наказав нам наш батько Йонадав.
JER|35|11|І сталося, коли Навуходоносор, цар вавилонський, прийшов був на цей Край, то ми сказали: Ходіть, і ввійдемо до Єрусалиму перед військом халдеїв та перед військом Араму. І осілися ми в Єрусалимі.
JER|35|12|І було слово Господа до Єремії таке:
JER|35|13|Так говорить Господь Саваот, Бог Ізраїлів: Іди, і скажеш до юдеянина та до мешканців Єрусалиму: Чи з цього не витягнете науки, щоб слухатися Моїх слів? говорить Господь.
JER|35|14|Додержано слова Єгонадава, Рехавового сина, що наказав був синам своїм не пити вина, і не пили вони аж до дня цього, бо послухалися наказу свого батька; а Я говорив до вас рано та пізно, та не слухалися ви Мене!
JER|35|15|І посилав Я до вас усіх Своїх рабів пророків рано та пізно, говорячи: Верніться но кожен зо своєї злої дороги, та виправте вчинки свої, і не ходіть за іншими богами, щоб служити їм, і сидіть на тій землі, що Я дав вам та вашим батькам! Та не схилили ви свого уха, і не послухались Мене.
JER|35|16|Бо додержали сини Єгонадава, сина Рехавового, наказа свого батька, що наказав був їм, а народ цей не послухався Мене.
JER|35|17|Тому так промовляє Господь Бог Саваот, Бог Ізраїлів: Ось Я спроваджую на Юду та на всіх мешканців Єрусалиму все те зло, що Я провіщав був про них. Бо Я говорив до них, та вони не слухали, і кликав Я їх, та вони не відповідали...
JER|35|18|А до дому Рехавітів Єремія сказав: Так говорить Господь Саваот, Бог Ізраїлів: За те, що ви слухалися наказа вашого батька Єгонадава, та держитеся всіх наказів його, і зробили те все, що Я заповів вам,
JER|35|19|тому так промовляє Господь Саваот, Бог Ізраїлів: Нема переводу в Йонадава, Рехавового сина, мужеві, що стоятиме перед лицем Моїм по всі дні!
JER|36|1|І сталося четвертого року Єгоякима, Йосіїного сина, царя Юдиного, було оце слово до Єремії від Господа, кажучи:
JER|36|2|Візьми собі книжкового звоя, і напиши на ньому всі ті слова, що Я говорив тобі про Ізраїля й про Юду, та про всі народи від дня, коли Я почав говорити тобі, від днів Йосії та аж до цього дня.
JER|36|3|Може почує дім Юдин усе те зло, що Я думаю вчинити їм, щоб вернулися кожен зо своєї злої дороги, а Я прощу їхню провину та їхній гріх.
JER|36|4|І покликав Єремія Баруха, Нерійїного сина, і Барух написав з уст Єремії всі Господні слова, що Він говорив йому, на книжковий звій.
JER|36|5|І наказав Єремія Барухові, кажучи: Я задержаний, не можу ввійти до Господнього дому.
JER|36|6|Тому піди сам, прочитай зо звою, що написав ти з моїх уст, Господні слова в вуха народу в Господньому домі в дні посту, а також в вуха всього Юди, що приходить зо своїх міст, відчитаєш їх.
JER|36|7|Може впаде їхнє благання перед Господнє лице, і вони вернуться кожен зо своєї злої дороги, бо великий гнів та лютість, що Господь говорив проти народу цього!
JER|36|8|І зробив Барух, син Нерійїн, усе, що наказав був йому пророк Єремія, щоб прочитати з книги Господні слова в Господньому домі.
JER|36|9|І сталося п'ятого року Єгоякима, Йосіїного сина, царя Юдиного, дев'ятого місяця, оголосили піст перед Господнім лицем для всього народу в Єрусалимі та для всього того народу, що поприходив з Юдиних міст до Єрусалиму.
JER|36|10|І прочитав Барух з книги Єреміїні слова в домі Господньому в кімнаті писаря Ґемарії, Шафанового сина, на горішньому подвір'ї, при вході до нової брами Господнього дому, в вуха всього народу.
JER|36|11|І почув Михей, син Ґемарії, Шафанового сина, всі Господні слова з книги,
JER|36|12|і зійшов до царського дому, до кімнати писаря, аж ось там сидять усі зверхники: писар Елішама, і Делая, син Шемаїн, і Елнатан, син Ахборів, і Ґемарія, син Шафанів, і Седекія, син Хананії, і всі зверхники.
JER|36|13|І розповів їм Михей всі ті слова, які він почув був, коли Барух читав із книги в вуха народу.
JER|36|14|І всі зверхники послали до Баруха Єгудія, сина Нетанії, сина Шелемії, сина Кушіїного, говорячи: Того звоя, що читав ти з нього в вуха народу, візьми його в свою руку та й прийди! І взяв Барух, син Нерійїн, звоя в свою руку та й прийшов до них.
JER|36|15|А ті сказали до нього: Сідай же, і прочитай його в наші вуха! І прочитав Барух в їхні вуха.
JER|36|16|І сталося, коли вони почули всі ці слова, жахнулися один перед одним, та й сказали Барухові: Конче перекажімо цареві всі ці слова!
JER|36|17|І запитали вони Баруха, говорячи: Розкажи нам, як ти писав усі ці слова з його уст?
JER|36|18|І сказав їм Барух: Він проказував мені з своїх уст усі ці слова, а я писав у книзі чорнилом.
JER|36|19|І сказали зверхники до Баруха: Іди, сховайся, ти та Єремія, і нехай ніхто не знає, де ви!
JER|36|20|І прийшли вони до царя на подвір'я, а звоя поклали в кімнаті писаря Елішами, і розповіли в вуха царя всі ті слова.
JER|36|21|І послав цар Єгудія взяти звоя, і той узяв його з кімнати писаря Елішами. І Єгудій прочитав його в вуха царя та в вуха всіх зверхників, що стояли при царі.
JER|36|22|А цар сидів у зимовому домі, дев'ятого місяця, і перед ним був розпалений коминок.
JER|36|23|І сталося, коли Єгудій перечитував три чи чотири стовпці, то цар відрізував це писарським ножем та й кидав до огню, що в коминку, аж поки не згорів увесь звій на огні, що в коминку...
JER|36|24|Та не злякалися й не роздерли своїх шат цар та всі його раби, що слухали всі ці слова.
JER|36|25|І хоч Елнатан, і Делая, і Ґемарія просили царя не палити того звою, та не послухався він їх.
JER|36|26|І наказав цар Єрахмеїлові, синові царевому, і Сераї, синові Азріїловому, і Шелемії, синові Авдіїловому, взяти писаря Баруха й пророка Єремію, та Господь їх сховав.
JER|36|27|І було Господнє слово до Єремії потому, як цар спалив був звоя та ті слова, що Барух написав з Єреміїних уст, говорячи:
JER|36|28|Візьми собі знову іншого звоя, і напиши на ньому всі перші слова, що були на першому звої, якого спалив Єгояким, цар Юдин.
JER|36|29|А про Єгоякима, царя Юдиного, скажеш: Так говорить Господь: Ти спалив цього звоя, говорячи: Нащо написав ти на ньому таке: Конче прийде цар вавилонський і знищить оцей Край, і вигубить в ньому людину й скотину.
JER|36|30|Тому так говорить Господь про Єгоякима, Юдиного царя: Не буде від нього сидячого на Давидовому троні, а його труп буде кинений на спекоту вдень та на холод вночі...
JER|36|31|І навіщу його та насіння його, і його рабів за їхні провини, і спроваджу на них та на мешканців Єрусалиму й на юдеянина все те зло, що Я говорив до них, та вони не послухали...
JER|36|32|І Єремія взяв іншого звоя, і дав його писареві Барухові, синові Нерійїному, і той написав на ньому з Єреміїних уст усі слова тієї книги, яку спалив був Єгояким, цар Юдин, в огні, і до них було додано ще багато подібних слів.
JER|37|1|І зацарював цар Седекія, син Йосійїн, замість Конії, сина Єгоякимового, якого зробив царем Навуходоносор, цар вавилонський, в Юдиному краї.
JER|37|2|Та не послухався ані він, ані його раби, ані народ Краю слів Господа, які Він говорив через пророка Єремію.
JER|37|3|І послав цар Седекія Єгухала, сина Шелеміїного, і священика Цефанію, сина Маасеїного, до пророка Єремії, говорячи: Помолися за нас до Господа, Бога нашого!
JER|37|4|А Єремія тоді ще вільно ходив серед народу, бо не дали його ще до в'язниці.
JER|37|5|А фараонове військо вийшло з Єгипту. І почули вістку про них халдеї, що облягали Єрусалим, і відійшли від Єрусалиму.
JER|37|6|І було слово Господнє до пророка Єремії, говорячи:
JER|37|7|Так промовив Господь, Бог Ізраїлів: Так скажете до Юдиного царя, що послав вас до мене поспитати мене: Ось фараонове військо, що вийшло вам на поміч, вернеться до свого краю, до Єгипту.
JER|37|8|А халдеї знову вернуться, і будуть воювати з цим містом, і здобудуть його, та й спалять його огнем.
JER|37|9|Так говорить Господь: Не обманюйте своїх душ, говорячи: Халдеї конче підуть від нас, бо не підуть вони.
JER|37|10|Бо якщо б ви побили все халдейське військо, що з вами воює, а з них залишилися б тільки ранені, то встане кожен із намету свого, і спалять це місто огнем...
JER|37|11|І сталося, коли халдейське військо відступило від Єрусалиму перед фараоновим військом,
JER|37|12|то вийшов Єремія з Єрусалиму, щоб піти до Веніяминового краю, і щоб сховатися там серед народу.
JER|37|13|Та коли він був біля Веніяминової брами, то був там начальник сторожі, а ім'я йому Їрійя, син Шелемеї, сина Хананіїного. І схопив він пророка Єремію, говорячи: Ти переходиш до халдеїв!
JER|37|14|А Єремія відказав: Неправда, я не переходжу до халдеїв! Та не послухав той його; і схопив Їрійя Єремію, і попровадив його до зверхників.
JER|37|15|І розгнівалися зверхники на Єремію, і побили його, та й віддали його до в'язниці в домі писаря Єгонатана, бо його зробили за в'язничний дім.
JER|37|16|І зійшов Єремія до темничної ями та до підвалу, і сидів там Єремія багато днів...
JER|37|17|І послав цар Седекія, і взяв його. І спитав його цар у своїм домі таємно й сказав: Чи є слово від Господа? І Єремія відказав: Є. І далі сказав: Ти будеш відданий в руку вавилонського царя...
JER|37|18|І сказав Єремія до царя Седекії: Що я згрішив тобі й рабам твоїм та цьому народові, що ви віддали мене до в'язниці?
JER|37|19|І де ваші пророки, що вам пророкували, говорячи: Цар вавилонський не прийде на вас та на Край цей?
JER|37|20|А тепер послухай, пане мій царю: хай упаде моє благання перед обличчя твоє, і не вертай мене до дому писаря Єгонатана, щоб не помер я там!...
JER|37|21|І наказав цар Седекія, й Єремію вмістили в подвір'ї в'язниці, і давали йому буханець хліба на день з вулиці пекарів, аж поки не скінчився ввесь хліб у місті. І сидів Єремія в подвір'ї в'язниці.
JER|38|1|І почув Шефатія, син Маттанів, і Ґедалія, син Пашхурів, і Юхал, син Шелемеїн, і Пашхур, син Малкійїн, ті слова, що Єремія говорив до всього народу, кажучи:
JER|38|2|Так говорить Господь: Хто сидітиме в цьому місті, той помре від меча, голоду та від моровиці, а хто вийде до халдеїв, той буде жити, і стане йому душа його за здобич, і він житиме!
JER|38|3|Так говорить Господь: Напевно буде дане це місто в руку війська вавилонського царя, і він здобуде його!
JER|38|4|І сказали зверхники до царя: Нехай же уб'ють цього чоловіка, бо він ослаблює руки вояків, позосталих у цьому місті, та руки всього народу, говорячи їм слова, як оці. Бо цей чоловік не шукає для цього народу добра, а тільки зла!...
JER|38|5|І сказав цар Седекія: Ось він у ваших руках, бо цар нічого не вдіє супроти вас.
JER|38|6|І взяли Єремію та й кинули його до ями Малкійї, царевого сина, що в подвір'ї в'язниці, і спустили Єремію шнурами. А в ямі була не вода, а тільки багно, і загруз Єремія в багні!
JER|38|7|І почув мурин Евед-Мелех, евнух, який був у царському домі, що Єремію кинули до ями, а цар сидів у Веніяминовій брамі.
JER|38|8|І вийшов Евед-Мелех з царського дому, та й сказав цареві, говорячи:
JER|38|9|Пане мій царю, ці люди вчинили зло в усьому, що зробили пророкові Єремії, якого кинули до ями, і помре він на своєму місці через голод, бо в місті нема вже хліба...
JER|38|10|І наказав цар муринові Евед-Мелехові, говорячи: Візьми з собою звідси троє люда, і витягнеш пророка Єремію з ями, поки він ще не вмер!
JER|38|11|І взяв Евед-Мелех тих людей з собою, і прийшов до царського дому під скарбницею, і набрав ізвідти подертого шмаття та непотрібних лахів, і спустив їх до Єремії до ями шнурами.
JER|38|12|І сказав мурин Евед-Мелех до Єремії: Поклади це подерте шмаття та лахи попід пахи своїх рук під шнури! І зробив Єремія так.
JER|38|13|І потягнули Єремію шнурами, і витягли його з ями. І сидів Єремія в подвір'ї в'язниці.
JER|38|14|І послав цар Седекія, і взяв пророка Єремію до себе, до третього входу, що в домі Господньому. І сказав цар до Єремії: Запитаю я тебе про щось, не заховуй від мене нічого!
JER|38|15|І сказав Єремія до Седекії: Коли я провіщу тобі, то чи справді не вб'єш ти мене? А коли пораджу тобі, то мене не послухаєш...
JER|38|16|І присягнув цар Седекія Єремії таємно, говорячи: Як живий Господь, що створив нам цю душу: не вб'ю тебе, і не дам тебе в руку тих людей, що шукають твоєї душі!
JER|38|17|І сказав Єремія до Седекії: Так говорить Господь, Бог Саваот, Бог Ізраїлів: Якщо справді вийдеш ти до зверхників вавилонського царя, то житиме душа твоя, а місто це не буде спалене огнем, і будеш жити ти та дім твій.
JER|38|18|А якщо ти не вийдеш до вавилонського царя, то це місто буде дане в руку халдеїв, і вони спалять його огнем, і ти не втечеш з їхньої руки...
JER|38|19|І сказав цар Седекія до Єремії: Я боюся юдеїв, що перейшли до халдеїв, щоб не дали мене в їхню руку, і щоб не насміялися з мене...
JER|38|20|І сказав Єремія: Не дадуть! Послухай Господнього голосу до того, що я говорю тобі, і буде добре тобі, і буде жити душа твоя!
JER|38|21|А якщо ти не схочеш вийти, то ось слово, що Господь мені виявив:
JER|38|22|І ось усі жінки, що залишилися в домі Юдиного царя, будуть відведені до зверхників вавилонського царя, і вони скажуть: Підмовили тебе й перемогли тебе твої приятелі; погрузили в багно твої ноги, та вони назад відійшли.
JER|38|23|А всі жінки твої та всі сини твої будуть відведені до халдеїв, і ти не втечеш з їхньої руки, бо рукою вавилонського царя будеш схоплений, а місто це буде спалене огнем...
JER|38|24|І сказав Седекія до Єремії: Нехай ніхто не знає про ці слова, і ти не помреш.
JER|38|25|Бо коли почують зверхники, що я говорив з тобою, то прийдуть до тебе та й скажуть тобі: Розкажи но нам, що говорив ти цареві! Не ховай перед нами, і не вб'ємо тебе. І що ж говорив тобі цар?
JER|38|26|то скажеш до них: Я склав своє благання перед царське обличчя, щоб не вертали мене до Єгонатанового дому, щоб там не померти.
JER|38|27|І прийшли всі зверхники до Єремії й запиталися його, і він розказав їм згідно зо всіма тими словами, що звелів був цар. І вони мовчки відійшли від нього, бо не довідались про обговорену річ.
JER|38|28|І сидів Єремія на подвір'ї в'язниці аж до дня, коли був здобутий Єрусалим. І сталося, як був здобутий Єрусалим:
JER|39|1|Дев'ятого року Седекії, царя Юдиного, місяця десятого, прийшов Навуходоносор, цар вавилонський, та все його військо до Єрусалиму та й облягли його.
JER|39|2|Одинадцятого року Седекії, місяця четвертого, дев'ятого дня місяця, був пробитий пролім до міста...
JER|39|3|І поприходили всі зверхники вавилонського царя, і посідали в Середущій брамі: Нерґал-Сар'ецер, Самгар, Нево, Сарсехім, старший евнух, Нерґал-Сар'ецер, старший маг, і вся решта зверхників вавилонського царя.
JER|39|4|І сталося, як побачив їх Седекія, цар Юдин, та всі вояки, то вони повтікали, і повиходили вночі з міста дорогою царського садка, брамою між обома мурами, і вийшли дорогою в степ.
JER|39|5|І погналося халдейське військо за ними, і догнали Седекію в єрихонських степах... І взяли вони його, і завели його до Навуходоносора, царя вавилонського, до Рівли, в краю Хамат, і той засудив його.
JER|39|6|І цар вавилонський порізав Седекіїних синів в Рівлі на очах його; і всіх шляхетних Юдиних порізав вавилонський цар...
JER|39|7|А очі Седекії він вибрав, і скував його мідяними кайданами, щоб відвести його до Вавилону...
JER|39|8|А дім царя та дому народу халдеї попалили огнем, і порозбивали мури Єрусалиму.
JER|39|9|А решту народу, позосталих у місті, та перебіжців, що попереходили до нього, і решту народу, що позосталися, вигнав Невузар'адан, начальник царської сторожі, до Вавилону.
JER|39|10|А з бідноти народу, що не мали нічого, Невузар'адан, начальник царської сторожі, позоставив декого в Юдиному краї, і дав їм того дня виноградники та поля.
JER|39|11|І наказав Навуходоносор, цар вавилонський, про Єремію, через начальника царської сторожі, говорячи:
JER|39|12|Візьми його, і зверни на нього свої очі, і не зроби йому нічого злого, і тільки як він скаже тобі, так з ним зроби!
JER|39|13|І послав Невузар'адан, начальник царської сторожі, і Невушазбан, старший евнух, і Нерґал-Сар'ецер, старший маг, та всі начальники вавилонського царя,
JER|39|14|і послали вони, і взяли Єремію з подвір'я в'язниці, і дали його до Ґедалії, сина Ахікама, сина Шафанового, щоб вивести його до дому. І осівся він серед народу.
JER|39|15|А до Єремії було Господнє слово, коли він був затриманий в подвір'ї в'язниці, таке:
JER|39|16|Іди, і скажеш до мурина Евед-Мелеха, говорячи: Так говорить Господь Саваот, Бог Ізраїлів: Ось Я наводжу Свої слова на це місто на зло, а не на добро, і вони будуть діятися перед тобою цього дня.
JER|39|17|Але тебе врятую цього дня, говорить Господь, і ти не будеш відданий в руку цих людей, яких ти боїшся.
JER|39|18|Бо конче врятую тебе, і від меча не впадеш ти, і буде тобі душа твоя за здобич, бо ти надіявся на Мене, говорить Господь.
JER|40|1|Слово, що було до Єремії від Господа по тому, як Невузар'адан, начальник царської сторожі, відпустив його з Рами, коли його він узяв, а він був закутий кайданами серед усього вигнання Єрусалиму та Юди, вигнаних до Вавилону.
JER|40|2|І взяв начальник царської сторожі Єремію, та й сказав до нього: Господь, Бог твій, говорив оце зло на це місце.
JER|40|3|І навів, і зробив Господь, як говорив був, бо ви згрішили Господеві, і не слухалися Його голосу, і сталася вам ця річ.
JER|40|4|А тепер ось я сьогодні розковую тебе з кайданів, що на твоїх руках. Якщо в очах твоїх добре піти зо мною до Вавилону, іди, і зверну я своє око на тебе. А якщо зле в твоїх очах піти зо мною до Вавилону, то залишись. Дивися, увесь Край перед тобою: куди тобі видається за добре й за справедливе піти, туди йди!
JER|40|5|І коли той не навертався на це, сказав далі: То вернися до Ґедалії, сина Ахікама, сина Шафанового, якого вчинив начальником вавилонський цар над Юдиними містами, і живи з ним серед народу; або куди тобі подобається, туди йди. І дав йому начальник царської сторожі їжі на дорогу та дарунка, і відпустив його.
JER|40|6|І прийшов Єремія до Ґедалії, сина Ахікамового, до Міцпи, й осівся з ним серед народу, позосталого в Краю.
JER|40|7|А коли всі військові зверхники, що були в полі, вони та їхні люди, прочули, що цар вавилонський учинив начальником над краєм Ґедалію, сина Ахікамового, і доручив йому мужчин і жінок та дітей, і тих з бідних Краю, що не були вигнані до Вавилону,
JER|40|8|то поприходили до Ґедалії до Міцпи: і Ізмаїл, син Нетаніїн, і Йоханан, та Йонатан, сини Кареахові, і Серая, син Танхуметів, і сини нетофеянина Ефая, і Єзанія, син маахеянина, вони та їхні люди.
JER|40|9|І Ґедалія, син Ахікама, сина Шафанового, заприсягнувся їм та їхнім людям, говорячи: Не бійтеся служити халдеям! Сидіть у Краї й служіть вавилонському цареві, і буде вам добре!
JER|40|10|А я ось сидітиму в Міцпі, щоб заступатися за вас перед халдеями, що прийдуть до нас. А ви збирайте вино й літні плоди та оливу, і складайте в ваш посуд, і сидіть у ваших містах, які ви зайняли!
JER|40|11|І також усі юдеї, що в Моаві й серед Аммонових синів, і в Едомі, і що в усіх краях, чули, що цар вавилонський полишив частину в Юді, і що вчинив над ними начальником Ґедалію, сина Ахікама, сина Шафанового.
JER|40|12|І вернулися всі юдеї зо всіх тих місць, куди були порозігнані, і прийшли до Юдиного краю, до Ґедалії до Міцпи, і зібрали вина та літніх плодів дуже багато.
JER|40|13|А Йоханан, син Кареахів, та всі військові зверхники, що були на полі, прийшли до Ґедалії до Міцпи,
JER|40|14|та й сказали до нього: Чи справді ти знаєш, що Бааліс, цар Аммонових синів, послав Ізмаїла, сина Нетаніїного, щоб убити тебе? Та не повірив їм Ґедалія, син Ахікамів.
JER|40|15|А Йоханан, син Кареахів, сказав таємно до Ґедалії в Міцпі, говорячи: Нехай я піду й уб'ю Ізмаїла, сина Нетаніїного, і ніхто про це не довідається. Нащо мають забити тебе, і буде розпорошений увесь Юда, зібраний до тебе, і погине останок Юди?
JER|40|16|І сказав Ґедалія, син Ахікамів, до Йоханана, сина Кареахового: Не роби цієї речі, бо лжу ти говориш на Ізмаїла!
JER|41|1|І сталося сьомого місяця, прийшов Ізмаїл, син Нетанії, сина Елішамового, з насіння царського, і вельможі царя, та десять люда з ним, до Ґедалії, Ахікамового сина, до Міцпи, і їли там разом хліб у Міцпі.
JER|41|2|І встав Ізмаїл, син Нетаніїн, і десять люда, що були з ним, та й ударили Ґедалію, сина Ахікама, сина Шафанового, мечем! І вбив він того, кого вавилонський цар настановив був начальником над Краєм...
JER|41|3|І повбивав Ізмаїл усіх юдеїв, що були з ним, з Ґедалією, у Міцпі, і халдеїв вояків, що знаходилися там.
JER|41|4|І сталося другого дня по вбивстві Ґедалії, а ніхто про це не знав,
JER|41|5|і поприходили люди з Сихему, з Шіло та з Самарії, вісімдесят люда оголенобородих, і в подертій одежі та з нарізаними знаками на тілі, а в їхній руці хлібна жертва та ладан, як принесення для Господнього дому.
JER|41|6|І вийшов Ізмаїл, син Нетаніїн, навпроти них з Міцпи, ідучи та плачучи. І сталося, коли він спіткав їх, то промовив до них: Прийдіть до Ґедалії, Ахікамового сина!
JER|41|7|І сталося, як прийшли вони до середини міста, то їх порізав Ізмаїл, син Нетаніїн, і повкидав їх до середини ями, він та ті люди, що були з ним...
JER|41|8|Та знайшлося між ними десять люда, і вони сказали до Ізмаїла: Не вбивай нас, бо ми маємо заховані в полі скарби: пшеницю, і ячмінь, і оливу, і мед. І той спинився, і не повбивав їх серед їхніх братів.
JER|41|9|А та яма, куди повкидав Ізмаїл усі трупи тих людей, була яма велика, яку зробив був цар Аса проти Баеші, Ізраїльського царя, її наповнив Ізмаїл, син Нетаніїн, трупами.
JER|41|10|І Ізмаїл узяв у полон усю решту народу, що був у Міцпі, царських дочок та ввесь народ, що зостався в Міцпі, якого Невузар'адан, начальник царської сторожі, доручив був Ґедалії, синові Ахікамовому. І забрав їх у полон Ізмаїл, син Нетаніїн, і пішов, щоб перейти до Аммонових синів.
JER|41|11|І почув Йоханан, син Кареахів, та всі військові зверхники, що були з ним, про все те зло, що зробив Ізмаїл, син Нетаніїн.
JER|41|12|І взяли вони всіх тих людей, і пішли воювати з Ізмаїлом, сином Нетаніїним, і знайшли його при великій воді, що в Ґів'оні.
JER|41|13|І сталося, як увесь народ, що був з Ізмаїлом, побачив Йоханана, сина Кареахового, та всіх військових зверхників, що були з ним, то зрадів.
JER|41|14|І відвернувся ввесь народ, якого взяв був до полону Ізмаїл з Міцпи, і вернулися, і пішли до Йоханана, сина Кареахового.
JER|41|15|А Ізмаїл, син Нетаніїн, утік з вісьмома людьми від Йоханана, і пішов до Аммонових синів.
JER|41|16|І взяв Йоханан, син Кареахів, та всі військові зверхники, що були з ним, усю решту народу, яку він вернув від Ізмаїла, сина Нетаніїного, з Міцпи, по тому, як той убив Ґедалію, сина Ахікамового, мужів вояків, і жінок, і дітей, і евнухів, що вернув з Ґів'ону.
JER|41|17|І пішли вони й стали на нічліг в Ґерут-Кімгамі, що при Віфлеємі, щоб піти й утікти до Єгипту
JER|41|18|від халдеїв, бо вони боялися їх, бо Ізмаїл, син Нетаніїв, убив Ґедалію, сина Ахікамового, якого вавилонський цар настановив був начальником над Краєм.
JER|42|1|І підійшли всі військові зверхники та Йоаханан, син Кареахів, і Єзанія, син Гошаїн, та ввесь народ від малого й аж до великого,
JER|42|2|та й сказали до пророка Єремії: Нехай упаде наше благання перед обличчя твоє, і молися за нас до Господа, Бога твого, за всю оцю решту, бо залишилося нас мало з багатьох, як бачать твої очі нас...
JER|42|3|І нехай виявить нам Господь, Бог твій, ту дорогу, якою ми підемо, та те діло, яке ми зробимо.
JER|42|4|І промовив до них пророк Єремія: Чую я! Ось я помолюся до Господа, вашого Бога, за вашими словами. І станеться, кожне слово, що Господь відповість вам, звіщу вам, нічого не затаю від вас.
JER|42|5|А вони сказали до Єремії: Нехай буде Господь проти нас за свідка правдивого та вірного, якщо ми не зробимо так, як усе те, з чим пошле тебе до нас Господь, Бог твій.
JER|42|6|Чи добре й чи зле, ми послухаємося голосу Господа, Бога нашого, що до Нього ми посилаємо тебе, щоб було нам добре, коли будемо слухатися голосу Господа, Бога нашого.
JER|42|7|І сталося з кінцем десятьох днів, і було Господнє слово до Єремії.
JER|42|8|І він покликав Йоханана, сина Кареахового, і всіх військових зверхників, що були з ним, та ввесь народ від малого й аж до великого,
JER|42|9|та й сказав до них: Так говорить Господь, Бог Ізраїлів, що ви послали мене до Нього скласти ваше благання перед Його лице:
JER|42|10|Якщо ви будете сидіти в цьому Краї, то збудую вас, а не розіб'ю, і засаджу вас, а не вирву, бо пожалував Я щодо того зла, що зробив був вам.
JER|42|11|Не бійтеся вавилонського царя, якого ви боїтеся, не бійтеся його, говорить Господь, бо з вами Я, щоб вас спасати, і щоб вас рятувати від його руки!
JER|42|12|І дам Я вам милість, і змилуюся над вами, і він верне вас до вашої землі.
JER|42|13|А якщо ви скажете: Не будемо сидіти в цьому Краї, щоб не слухатися голосу Господа, Бога вашого,
JER|42|14|кажучи: Ні, ми підемо до єгипетського краю, де не побачимо війни, і не почуємо звуку сурми, і на хліб не будемо голодні, і там будемо сидіти,
JER|42|15|то тому послухайте тепер Господнього слова, решто Юдина! Так говорить Господь Саваот, Бог Ізраїлів: Якщо ви справді скеруєте своє обличчя, щоб іти до Єгипту, і ввійдете, щоб чужинцями замешкати там,
JER|42|16|то станеться: той меч, що ви боїтеся його, досягне вас там, ув єгипетськім краї, а голод, якого ви лякаєтесь, пристане до вас в Єгипті, і там ви повмираєте...
JER|42|17|І станеться, всі люди, що звернули своє обличчя на мандрівку до Єгипту, щоб чужинцями замешкати там, повмирають від меча, від голоду та від моровиці, і жоден з них не позостанеться й не втече через те зло, що Я спроваджу на них...
JER|42|18|Бо так каже Господь, Саваот, Бог Ізраїлів: Як вилився гнів Мій та лютість Моя на мешканців Єрусалиму, так виллється лютість Моя на вас, коли ви прийдете до Єгипту, і будете там на клятьбу, і на застрашення, і на прокляття, і на ганьбу, і ви вже не побачите цього місця...
JER|42|19|Господь говорить до вас, Юдина решто: Не ходіть до Єгипту! Добре знайте, що сьогодні Я вас остеріг!
JER|42|20|Бо ви зблудилися в душах своїх, що послали мене до Господа, вашого Бога, говорячи: Молися за нас до Господа, Бога нашого, і все, що скаже Господь, Бог наш, так перекажи нам, і ми зробимо.
JER|42|21|І переказав я вам сьогодні, та не послухалися ви голосу Господа, Бога вашого, та всього того, з чим послав Він мене до вас.
JER|42|22|А тепер знайте напевно, що повмираєте від меча, голоду та від зарази в тому місці, куди хочете йти, щоб жити там чужинцями...
JER|43|1|І сталося, як Єремія скінчив говорити до всього народу всі слова Господа, Бога їхнього, всі ті слова, з якими послав його до них Господь, Бог їхній,
JER|43|2|то сказав Азарія, син Гошаїн, і Йоханан, син Кареахів, та всі бундючні люди, кажучи до Єремії: Брехню ти говориш! Не послав тебе Господь, Бог наш, сказати: Не входьте до Єгипту, щоб чужинцями замешкати там,
JER|43|3|то тебе намовив проти нас Барух, син Нерійїн, щоб віддати нас у руку халдеїв, щоб повбивати нас, і щоб вигнати нас до Вавилону...
JER|43|4|І не послухався Йоханан, син Кареахів, і всі військові зверхники та ввесь народ Господнього голосу, щоб сидіти в Юдиному краї.
JER|43|5|І взяв Йоханан, син Кареахів, та всі військові зверхники всю Юдину решту, що вернулися від усіх народів, куди були вигнані, щоб замешкати в Юдиному краї,
JER|43|6|мужчин та жінок, і дітей та царських дочок, і всяку душу, що Невузар'адан, начальник царської сторожі, позоставив був із Ґедалією, сином Ахікама, сина Шафанового, і з пророком Єремією та з Барухом, сином Нерійїним,
JER|43|7|і прийшли до єгипетського краю, бо не послухалися Господнього голосу, і прийшли до Тахпанхесу.
JER|43|8|І було слово Господнє до Єремії в Тахпанхесі таке:
JER|43|9|Візьми в свою руку великі каміння, і сховай їх у глині на цегляному майдані, що при вході до фараонового дому в Тахпанхесі, на очах юдейських людей.
JER|43|10|І скажеш до них: Так говорить Господь Саваот, Бог Ізраїлів: Ось Я пошлю й візьму Навуходоносора, царя вавилонського, Мого раба, і поставлю його трона над тими каміннями, що Я поховав, і він своє царське шатро розтягне над ними.
JER|43|11|І він прийде, і вдарить єгипетський край: що призначене на смерть піде на смерть, а що до полону до полону, а що на меча піде на меча...
JER|43|12|І підпалю огонь у домах єгипетських богів, і він попалить їх, і забере їх у полон, і він очистить єгипетський край, як чистить пастух свою одіж, і вийде звідти в спокої...
JER|43|13|І він поламає посвячені стовпи Бет-Шемеша, що в єгипетському краї, а доми єгипетських богів попалить огнем.
JER|44|1|Слово, що було до Єремії про всіх юдеїв, що сиділи в єгипетському краї, що сиділи в Міґдолі, і в Тахпанхесі, і в Нофі, і в краю Патрос, говорячи:
JER|44|2|Так говорить Господь Саваот, Бог Ізраїлів: Ви бачили все те зло, що Я спровадив на Єрусалим та на всі Юдині міста, і ось вони цього дня руїна, і немає в них мешканця...
JER|44|3|Це через їхнє зло, яке вони зробили, щоб гнівити Мене, ходячи кадити, служити іншим богам, яких не знали ані вони, ані ви, ані ваші батьки.
JER|44|4|І посилав Я до вас усіх Моїх рабів пророків, рано та пізно, кажучи: Не робіть цієї обридливої речі, яку Я зненавидив!
JER|44|5|Та не слухали вони, і не нахилили уха свого, щоб відвернутися від свого зла, щоб не кадити іншим богам.
JER|44|6|І вилилась лютість Моя та Мій гнів, і запалав він в Юдиних містах та на вулицях Єрусалиму, і стали вони руїною та пустинею, як бачите цього дня...
JER|44|7|А тепер так говорить Господь, Бог Саваот, Бог Ізраїлів: Нащо ви робите велике зло своїм душам, вигублюючи собі чоловіка та жінку, дитину й немовля з-серед Юди, щоб не залишилася вам решта?
JER|44|8|Нащо ви робите, щоб гнівити Мене чинами рук своїх, щоб кадити іншим богам в єгипетському краї, куди ви прийшли чужинцями замешкати там, щоб погубити себе, і щоб стати прокляттям та ганьбою серед усіх людів землі?
JER|44|9|Чи забули ви зло ваших батьків, та зло Юдиних царів, і зло жінок його, і зло ваше та зло ваших жінок, що наробили в Юдиному краї та на вулицях Єрусалиму?
JER|44|10|Не були вони впокорені аж до цього дня, і не бояться, і не ходять Законом Моїм та Моїми уставами, що Я дав вам та вашим батькам.
JER|44|11|Тому так промовляє Господь Саваот, Бог Ізраїлів: Ось Я зверну обличчя Своє на вас вам на зло, щоб викоренити всього Юду!
JER|44|12|І візьму Я залишок Юди, що звернули обличчя своє на мандрівку в єгипетський край, щоб чужинцями замешкати там, і погинуть усі в єгипетському краї, попадають від меча та від голоду, погинуть від малого й аж до великого, повмирають від меча та від голоду, і стануть клятьбою, застрашенням, і прокляттям та ганьбою...
JER|44|13|І покараю замешкалих в єгипетському краї, як покарав Я Єрусалим, мечем, голодом та моровицею...
JER|44|14|І не буде втікача та врятованих із решти Юди, що прийшли чужинцями замешкати там в єгипетському краї, щоб вернутися до Юдиного краю, куди вони бажають усією душею своєю вернутися й оселитися там. Але не вернуться вони, хіба тільки поодинокі втікачі!
JER|44|15|І відповіли Єремії всі ті люди, що знали, що їхні жінки кадять іншим богам, і всі ті жінки, що стояли там, великий збір, і ввесь народ, що сидів в єгипетському краї в Патросі, говорячи:
JER|44|16|Щодо слова, що ти говорив до нас Господнім Ім'ям, ми не слухаємо тебе.
JER|44|17|Бо напевно виконаємо кожне те слово, що виходить із наших уст, щоб кадити небесній цариці й лити їй литі жертви, як робили ми та батьки наші, царі наші та зверхники наші в Юдиних містах та на вулицях Єрусалиму. І насичувалися ми хлібом, і було нам добре, а зла ми не бачили.
JER|44|18|А відколи перестали ми кадити небесній цариці й лити ій литі жертви, брак нам усього, і ми гинемо від меча та голоду!
JER|44|19|А коли ми кадимо небесній цариці й приносимо їй литі жертви, то хіба без відома наших чоловіків ми робимо для неї жертовні калачі з її зображенням, і ллємо їй литі жертви?
JER|44|20|І сказав Єремія до всього народу, до чоловіків та до жінок, та до всього народу, що відповідали йому таке, говорячи:
JER|44|21|Хіба не кадило, яке кадили в Юдиних містах та на вулицях Єрусалиму ви та ваші батьки, ваші царі та зверхники ваші й народ цього краю, хіба не згадав це Господь, і не ввійшло воно до серця Його?
JER|44|22|І не зміг Господь більше знести зла ваших чинів, та ті гидоти, що ви наробили, тому став ваш Край руїною, і застрашенням та прокляттям, так що немає мешканця, як бачите цього дня...
JER|44|23|За те, що кадили ви, і що грішили Господеві, і не слухалися Господнього голосу, і не ходили Законом Його й Його правом та свідоцтвами Його, тому спіткало вас оце зло, як бачите цього дня.
JER|44|24|І сказав Єремія до всього народу та до всіх жінок: Послухайте Господнього слова, ввесь Юдо, що в єгипетському краї!
JER|44|25|Так говорить Господь Саваот, Бог Ізраїлів, кажучи: Ви та ваші жінки говорили своїми устами й своїми руками виконували, кажучи: Конче виконаємо свої присяги, що ми присягали кадити небесній цариці й лити їй литі жертви, тому напевно здійсніте ваші присяги, і конче виконайте обітниці ваші.
JER|44|26|Тому то послухайте Господнього слова, ввесь Юдо, що сидиш в єгипетському краї: Ось Я присягнув великим Своїм Ім'ям, говорить Господь, що не буде вже Ім'я Моє кликатися устами жодного юдеянина, кажучи: Живий Господь Бог! у всьому єгипетському краї.
JER|44|27|Ось Я пильную вас на зло, а не на добро, і загине кожен юдеянин, що в єгипетському краї, від меча та від голоду, аж до їх скону.
JER|44|28|А врятовані від меча вернуться з єгипетського краю до краю Юдиного нечисленними. І пізнає ввесь останок Юди, що прийшли до єгипетського краю чужинцями замешкати там, чиє слово виконається: Моє чи їхнє?
JER|44|29|А оце вам той знак, говорить Господь, що Я відвідаю вас у цьому місці, щоб ви пізнали, що конче справдяться Мої слова на вас на зло.
JER|44|30|Так говорить Господь: Ось Я видам фараона Хофру, єгипетського царя, в руку його ворогів та в руку тих, що шукають душі його, як дав Я Седекію, Юдиного царя, у руку Навуходоносора, вавилонського царя, його ворога, що шукав душі його!
JER|45|1|Слово, що говорив пророк Єремія до Баруха, Нерійїного сина, коли той писав ці слова в книзі з Єреміїних уст, за четвертого року Єгоякима, сина Йосіїного, царя Юдиного, кажучи:
JER|45|2|Так говорить Господь, Бог Ізраїлів, про тебе, Баруху:
JER|45|3|Ти сказав був: Ой горе мені, бо додав Господь смутку до болю мого! Я змучивсь зідханням своїм, і не знайшов відпочинку!
JER|45|4|Так скажеш йому: Так говорить Господь: Ось Я поруйную, що Я збудував, а що Я насадив, те Я вирву, також усю землю Свою.
JER|45|5|А ти ось шукаєш для себе великого. Не шукай, бо ось Я наведу зло на кожне тіло, говорить Господь, а тобі дам душу твою за здобич на всіх тих місцях, де ти будеш ходити!
JER|46|1|Слово Господнє, що було пророкові Єремії про народи.
JER|46|2|На Єгипет. На військо фараона Нехо, єгипетського царя, що був над річкою Ефратом у Каркеміші, якого побив Навуходоносор, вавилонський цар, за четвертого року Єгоякима, сина Йосіїного, царя Юдиного:
JER|46|3|Приготуйте щитка та щита, і приступіть до війни!
JER|46|4|Запрягайте но коні й сідайте, верхівці, і поставайте в шоломах! Вичистіть ратища та зодягніться в кольчуги!
JER|46|5|Що то бачу: вони полякались й назад відступають? А лицарі їхні подолані та втікають і не оглядаються... Страхіття навколо, говорить Господь!
JER|46|6|Швидкий не втече, і не врятується лицар, на півночі, при річці Ефраті спіткнуться вони та й попадають!
JER|46|7|Хто то такий підіймається, мов та Ріка, як річки, його води хвилюються?
JER|46|8|Єгипет, немов та Ріка, підіймається він, мов річки, його води хвилюються, і каже: Підіймуся, покрию я землю, і вигублю місто й мешканців його!
JER|46|9|Сідайте на коні й шалійте, колесниці! І хай лицарі вийдуть, Куш та Пут, що хапають щита, та людійці, що хапають, натягують лука!
JER|46|10|А день цей Господа, Бога Саваота, день помсти, щоб помститися над ворогами Своїми, і меч буде жерти й насититься, і досить нап'ється їхньої крови, бо це буде жертва для Господа, Бога Саваота, в північному краї при річці Ефраті!
JER|46|11|Піди до Ґілеаду, й бальзаму візьми, дівчино, дочко Єгипту! Надармо вживаєш ти ліків багато, своїх ран не загоїш!
JER|46|12|Почули народи про ганьбу твою, а крику твого стала повна земля, бо спіткнулися лицар об лицаря, разом упали обоє вони!
JER|46|13|Слово, що говорив Господь пророкові Єремії про прихід Навуходоносора, царя вавилонського, щоб побити єгипетську землю:
JER|46|14|Розкажіте в Єгипті, і розголосіте в Міґдолі, і розголосіте в Нофі й Тахпанхесі! Скажіть: стань, і собі приготуйся, бо меч пожирає круг тебе!
JER|46|15|Чому твої лицарі впали? Не втрималися, бо пхнув їх Господь!...
JER|46|16|Стало багато таких, що спіткнулися, навіть падають один на одного й говорять: Уставай, і до свого народу вернімось, і до краю народження нашого, перед згубним мечем!
JER|46|17|Назвіте ім'я фараону, цареві єгипетському: Загибіль, пропустив він усталений час!
JER|46|18|Як живий Я, каже Цар, що Господь Саваот Йому Ймення, він прийде, немов би Фавор у горах, й як при морі Кармел!
JER|46|19|Приготуй необхідне собі на мандрівки, мешканко, о дочко Єгипту, бо стане спустошенням Ноф, і він спалений буде, і в ньому не буде мешканця!
JER|46|20|Єгипет теля гарноусте, та летить он із півночі ґедзь!...
JER|46|21|Серед нього й його наймити, мов телята вгодовані, та й вони повернулись назад, повтікали разом, не спинились, бо день їхнього нещастя прийшов ось на них, час навіщення їх...
JER|46|22|Розлягається голос його, як гадюче сичання, бо йдуть вони з військом, і прийдуть до нього з сокирами, мов дроворуби...
JER|46|23|Вони ліс його витнуть, говорить Господь, хоч він непрохідний, бо стануть вони більш численні, як та сарана, і не буде числа їм.
JER|46|24|Засоромлена буде єгипетська донька, буде видана в руку народу північного...
JER|46|25|Говорить Господь Саваот, Бог Ізраїлів: Ось Я покараю Амона із Но, і фараона, і Єгипет, і богів його, і царів його, і фараона, і тих, що на нього надіються.
JER|46|26|І дам їх у руку всіх тих, хто шукає їхню душу, і в руку Навуходоносора, царя вавилонського, і в руку рабів його, а потому він буде заселений, як за днів давніх, говорить Господь!
JER|46|27|А ти не лякайся, рабе Мій Якове, і не страшися, Ізраїлю, бо Я ось врятую тебе здалека, і насіння твоє з краю їхнього полону! І вернеться Яків, і буде спокійний, і буде безпечний, і не буде того, хто б його настрашив!
JER|46|28|А ти не лякайся, рабе Мій Якове, каже Господь, бо Я з тобою, бо зроблю Я кінець всім народам, куди тебе вигнав, та з тобою кінця не зроблю, і тебе покараю за правом, і тебе непокараним не полишу!
JER|47|1|Слово Господнє, що було пророкові Єремії на филистимлян, перше як фараон побив Аззу.
JER|47|2|Так говорить Господь: Ось підіймаються води із півночі, і стануть вони за потік заливний, і заллють вони землю та все, що на ній, місто й замешкалих в ньому, і буде кричати людина, і кожен мешканець землі заголосить...
JER|47|3|Через гук тупотіння копит баских коней його, через гуркіт його колесниць, через скрип його кіл не звернулись батьки до синів, бо зомліли їм руки,
JER|47|4|бо настав це той день, щоб понищити всіх филистимлян, щоб Тиру й Сидонові вигубити помічну всяку рештку... Бо понищить Господь филистимлян, рештку острова Кафтора,
JER|47|5|шолудивою стане Азза, згине Ашкелон, решта долини їхньої... Як довго ти будеш нарізи робити собі у жалобі?
JER|47|6|О мечу Господній, аж доки ти не заспокоїшся? Вернися до піхви своєї, заспокойся й замовкни!
JER|47|7|Але як заспокоїться він, коли наказав йому це Сам Господь? До Ашкелону й до берегу моря, туди Він призначив його!...
JER|48|1|На Моава. Так каже Господь Саваот, Бог Ізраїлів: Горе місту Нево, бо воно поруйноване; Кір'ятаїм посоромлений, здобутий; посоромлений Замок високий, заляканий...
JER|48|2|Нема більше слави Моаву! У Хешбоні лихе вимишляють на нього: Ходімо, і витнім його із народу! Теж, Мадмене, замовкнеш і ти: за тобою йде меч!
JER|48|3|Чути крик із Горонаїму: Руїна й нещастя велике!
JER|48|4|Моав поруйнований, крик підняли аж до Цоару,
JER|48|5|бо ходом в Лухіт підуть догори з великим плачем, бо на збіччі Горонаїму чути крик боязкий про руїну...
JER|48|6|Утікайте, рятуйте хоч душу свою, і станете, мов отой верес в пустині!
JER|48|7|Бо за те, що надіявся ти на вчинки свої та на скарби свої, ти також будеш узятий, і піде Кемош до полону, а разом із ним його священики та його зверхники...
JER|48|8|І прийде руїна до кожного міста, і не буде врятоване жодне із них, і загине долина, й погублена буде рівнина, бо так говорив був Господь!...
JER|48|9|Дайте крила Моаву, і він відлетить, і міста його стануть спустошенням, так що не буде мешканця у них...
JER|48|10|Проклятий, хто робить роботу Господню недбало, і проклятий, хто від крови на меча свого стримує!
JER|48|11|Спокійний Моав від юнацтва свого, і мирний на дріжджах своїх, і не лито із посуду в посуд його, і він на вигнання не йшов, тому в нім його смак позостався, а запах його не змінився.
JER|48|12|Тому то ось дні настають, говорить Господь, і пошлю Я на нього розливачів, і його розіллють, і посуд його опорожнять, і дзбанки його порозбивають!...
JER|48|13|І за Кемоша Моав посоромлений буде, як Ізраїлів дім посоромлений був за Бет-Ел, за місце надії своєї.
JER|48|14|Як говорите ви: Ми хоробрі та сильні до бою?
JER|48|15|Попустошений буде Моав, і до міст його ворог підійметься, і підуть добірні його юнаки на заріз, каже Цар, що Господь Саваот Йому Ймення...
JER|48|16|Близький похід нещастя Моава, а лихо його дуже квапиться...
JER|48|17|Співчувайте йому, всі довкілля його, і всі, хто ім'я його знає, скажіть: Як зламалося сильне це берло, ця палиця пишна!
JER|48|18|Спустися зо слави своєї, і всядься в пустині, о мешканко, дочко Дівону, бо спустошник Моава до тебе прийшов, і понищив твердині твої!
JER|48|19|Стань на дорозі й чекай, мешканко Ароеру, питай втікача та врятовану, кажи: Що це сталося?
JER|48|20|Моав посоромлений, бо розтрощений він, ридайте та плачте, і звістіте в Арноні, що Моав попустошений!
JER|48|21|І суд ось прийшов на рівнинний цей край, на Холон й на Ягцу, і на Мефаат,
JER|48|22|і на Дівон, і на Нево, і на Бет-Дівдатаїм,
JER|48|23|і на Кір'ятаїм, і на Бет-Ґамул, і на Бет-Меон,
JER|48|24|і на Керіййот, і на Боцру, і на всі міста моавського краю, далекі й близькі...
JER|48|25|І відтятий Моавові ріг, і рамено його розтрощене, говорить Господь.
JER|48|26|Упійте його, бо пишавсь проти Господа він, і він з плюскотом упаде до блювоти своєї, і станеться й він посміховиськом!...
JER|48|27|І чи ж для тебе Ізраїль не був посміховиськом цим? Хіба серед злодіїв був знайдений він, що ти скільки говориш про нього, то все головою хитаєш?
JER|48|28|Покиньте міста, й пробувайте на скелі, мешканці Моава, і будьте, немов та голубка, що над краєм безодні гніздиться!
JER|48|29|Ми чули про гордість Моава, що чванливий він дуже, про надутість його і його гордування, про бундючність його та пиху його серця.
JER|48|30|Я знаю, говорить Господь, про зухвальство його, і про його балачки безпідставні, робили вони неслухняне!
JER|48|31|Ридаю тому над Моавом, і кричу за Моавом усім, зідхаю над людьми Кір-Хересу...
JER|48|32|Більш як за Язером Я плакав, Я плакатиму за тобою, винограднику Сівми! Галузки твої перейшли аж за море, досягли аж до моря Язера. Спустошник напав на осінній твій плід, і на винобрання твоє,
JER|48|33|і забрана буде потіха твоя та радість твоя з виноградника й з краю Моава, і вино із чавила спиню! Не буде топтати топтач, радісний крик при збиранні не буде вже радісним криком збирання...
JER|48|34|Від крику Хешбону аж до Ел'але, аж до Ягацу нестися буде їхній голос, від Цоару аж до Горонаїму, до Еґлат-Шелішійї, бо й вода із Німріму пустинею стане...
JER|48|35|І вигублю Я із Моава, говорить Господь, того, хто для жертов виходить на пагірок, і богові кадить своєму.
JER|48|36|Тому стогне серце Моє за Моавом, немов та сопілка, і стогне серце Моє, як сопілка, за людьми Кір-Хересу, бо погинули ті, хто багатство набув!...
JER|48|37|Тому кожна голова облисіла, і кожна борода обстрижена, на руках у всіх порізи жалоби, і на стегнах верета...
JER|48|38|На всіх дахах Моава й на площах його самий лемент, бо розбив Я Моава, мов посуд, якого не люблять, говорить Господь...
JER|48|39|Як він розтощений плачуть, як ганебно Моав утікав, і як він посоромлений! І Моав став за посміх та пострах для всього довкілля його!
JER|48|40|Бо так промовляє Господь: Ось він, як орел, прилетить, і крила свої над Моавом розгорне,
JER|48|41|міста будуть взяті, й твердині захоплені... І того дня стане серце лицарства Моава, як серце жони-породіллі!
JER|48|42|І з народів Моав буде вигублений, бо пишавсь проти Господа він...
JER|48|43|Страх, та безодня, та пастка на тебе, мешканче Моава! говорить Господь.
JER|48|44|Хто від страху втече, той в безодню впаде, хто ж з безодні підійметься, той буде схоплений в пастку... Бо спроваджу на нього, на того Моава, рік їхньої кари, говорить Господь.
JER|48|45|Втікачі знесилені будуть ставати у тіні Хешбону, бо вийде огонь із Хешбону, а полум'я з-поміж Сигону, і поїсть край волосся на скроні Моаву та череп синів галасливих...
JER|48|46|Горе, Моаве, тобі! Загинув Кемошів народ, бо сини твої взяті в полон, твої ж дочки в неволю!...
JER|48|47|І верну Я Моавові долю наприкінці днів, говорить Господь. Аж досі суд на Моава.
JER|49|1|На Аммонових синів. Так говорить Господь: Чи немає синів у Ізраїля? Чи немає спадкоємця в нього? Чому Ґада Мілком одідичив й осівся народ його по містах його?
JER|49|2|Тому настають ось дні, говорить Господь, і Я розголошу крик військовий на Раббу Аммонових синів, і вона стане за купу руїн, а підлеглі міста її спалені будуть огнем, і знов одідичить Ізраїль спадок свій, говорить Господь.
JER|49|3|Ридай, о Хешбоне, бо місто зруйноване! Кричіть, дочки Рабби, опережіться веретою, лементуйте й блукайте по обійстях, бо Мілком до полону іде, його священики й його зверхники разом!
JER|49|4|Чого ти долинами хвалишся? Долина твоя розпливається кров'ю, о дочко невірна, що на скарби свої покладаєш надію та кажеш: Хто прийде до мене?
JER|49|5|Ось Я страх припроваджу на тебе, говорить Господь, Бог Саваот, із усього довкілля твого, і ви повтікаєте кожен наперед себе, і не буде кому втікачів позбирати!...
JER|49|6|А потім верну Я долю Аммонових синів, говорить Господь.
JER|49|7|На Едома. Так говорить Господь Саваот: Чи в Темані немає вже мудрости? Чи згинула рада розумних? Хіба зіпсувалась їхня мудрість?
JER|49|8|Утікайте, оберніться плечима, сядьте глибше, мешканці Дедану, бо привів Я нещастя Ісава на нього, той час, коли покараю його!
JER|49|9|Якщо прийдуть до тебе збирачі винограду, вони не полишать останків, якщо ж прийдуть злодії вночі, напсують, скільки схочуть.
JER|49|10|Бо обнажив Я Ісава, повідкривав усі криївки його, і він сховатись не зможе, спустошене буде насіння його, й його браття, і сусіди його, і не буде його!
JER|49|11|Залиши свої сироти, Я утримаю їх при житті, а вдови твої хай надію на Мене кладуть!
JER|49|12|Бо так промовляє Господь: Ось і ті, що не мали б пити чаші цієї, пити будуть напевне, а ти непокараним будеш? Не будеш без кари, бо справді ти питимеш чашу!
JER|49|13|Бо Собою присяг Я, говорить Господь, що Боцра за спустошення стане, за ганьбу, пустиню й прокляття, і руїнами вічними стануть міста її всі!
JER|49|14|Я звістку від Господа чув, і відправлений вісник між люди: Зберіться й прийдіть проти неї, і встаньте на бій,
JER|49|15|бо тебе Я зробив ось малим між народами, погордженим серед людей!
JER|49|16|Страхіття твоє обманило тебе й гордість серця твого, тебе, що в розщілинах скелі живеш, що високих підгірків тримаєшся. Та коли б ти кубло своє й високо звив, мов орел, то й ізвідти Я скину тебе, промовляє Господь.
JER|49|17|І стане Едом за страхіття, кожен, хто буде проходити ним, остовпіє й засвище, як порази його всі побачить...
JER|49|18|Як Содом та Гоморру й сусідів її поруйновано, каже Господь, так ніхто там не буде сидіти, і не буде в нім мешкати чужинцем син людський.
JER|49|19|Ось підійметься він, немов лев, із темного лісу Йордану на водяні луки, і Я вмент зроблю, що він побіжить геть від них, а хто вибраний буде, того Я поставлю над ними. Бо хто є подібний Мені, і хто покличе Мене перед суд, і хто пастир такий, що перед обличчям Моїм устоїть?
JER|49|20|Тому то послухайте задум Господній, що Він на Едома задумав, і думки Його ті, які Він на мешканців Теману замислив: Направду, найменших з отари потягнуть, і попустошать пасовисько їхнє при них!
JER|49|21|Від гуку упадку їхнього буде тремтіти земля, буде зойк, аж на морі Червоному чути їхній голос.
JER|49|22|Ось підійметься він, як орел, і літатиме, й крила свої над Боцрою розгорне: і стане серце хоробрих едомлян в той день, немов серце жони-породіллі...
JER|49|23|На Дамаск. Засоромивсь Хамаш та Арпад, бо злу звістку почули; в неспокої тривожнім вони, як те море, що не може вспокоїтись.
JER|49|24|Дамаск сторопів, обернувся втікати, і страх його міцно охопив, біль та муки його обгорнули, немов породіллю...
JER|49|25|Як спорожніло славне це місто, місто втіхи Моєї!
JER|49|26|Тому юнаки його падати будуть на площах його, і всі військові погинуть того дня, говорить Господь Саваот.
JER|49|27|І під муром Дамаску огонь запалю, і він пожере Бен-Гададські палаци!...
JER|49|28|На Кедар та на царства Хацору, що їх побив Навуходоносор, цар вавилонський. Так говорить Господь: Уставайте, ідіть на Кедар, і нехай попустошать війська синів сходу!
JER|49|29|Заберуть їхні намети та їхню отару, їхні покрови та всі їхні речі, та їхніх верблюдів собі заберуть, і над ними кричатимуть: Жах звідусіль!
JER|49|30|Утікайте, мандруйте скоріш, сховайтесь в глибоке, мешканці Хацору, говорить Господь, бо раду нарадив на вас Навуходоносор, цар вавилонський, і задум задумав на вас!
JER|49|31|Уставайте, ідіть на народ, що спокійно, безпечно живе, промовляє Господь, немає воріт, і нема в нього засувів, самітно живуть.
JER|49|32|І стануть верблюди їхні здобиччю, а їхні череда грабежем, і на всі вітри розвію Я їх, хто волосся довкола стриже, і зо всіх їхніх сторін припроваджу на них їхню погибіль, говорить Господь...
JER|49|33|І стане Хацор за мешкання шакалів, за вічне спустошення, не замешкає там людина, і син людський не спиниться в ньому!...
JER|49|34|Слово Господнє, що було пророкові Єремії на Елам на початку царювання Седекії, Юдиного царя, таке:
JER|49|35|Так говорить Господь Саваот: Ось Я зламаю еламського лука, головну їхню силу!
JER|49|36|І з чотирьох кінців неба спроваджу чотири вітри до Еламу, і їх розпорошу на всі ці вітри, і не буде такого народу, куди б не прийшли ці вигнанці з Еламу...
JER|49|37|І настрашу Елам перед їхніми ворогами та перед всіма, хто їхню душу шукає, і лихо на них наведу, лютість гніву Мого, говорить Господь, і пошлю Я за ними меча, аж поки не вигублю їх!
JER|49|38|І поставлю Престола Свого в Еламі, і вигублю звідти царя й його зверхників, каже Господь...
JER|49|39|Але буде наприкінці днів, поверну Я Еламові долю, говорить Господь.
JER|50|1|Слово, що Господь говорив на Вавилон, на землю халдеїв через пророка Єремію:
JER|50|2|Звістіть між народами й розголосіть, підійміте прапора та розголосіть, не затайте, скажіть: Здобутий уже Вавилон, засоромлений Бел, зламаний Меродах, боввани його посоромлені, порозбивані всі його божища!
JER|50|3|Бо на нього із півночі вийшов народ, що оберне в спустошення землю його, і не буде мешканця у нім: від людини та аж до скотини, усі помандрують та підуть!...
JER|50|4|За тих днів і того часу, говорить Господь, поприходять сини Ізраїлеві, разом вони й сини Юди, усе плачучи, будуть ходити та Господа, Бога свого шукати...
JER|50|5|Вони будуть питати про Сіона, куди їхні обличчя повернені, щоб прийти й прилучитись до Господа вічним заповітом, який не забудеться!
JER|50|6|Мій народ це отара загинула: пастирі їхні вчинили блудячими їх, їх загнали на гори, й ходили вони від гори до підгір'я, забули про ложе своє...
JER|50|7|Усі, що знаходили їх, жерли їх, і противники їхні говорили: Не завинимо за те, бо вони прогрішилися Господу, Пасовиську правди й надії батьків їхніх, Господеві.
JER|50|8|Біжіть з Вавилону, і виходьте із краю халдеїв, і будьте, як козлята ті перед отарою!
JER|50|9|Бо ось Я позбуджую, і на Вавилон наведу збір великих народів з північного краю, і вони проти нього шикуються, звідти здобутий він буде! Його стріли, мов лицар, якому щастить, не вертаються дармо,
JER|50|10|і здобиччю стане Халдея, наситяться всі, хто пустошить її, промовляє Господь...
JER|50|11|Бо радієте ви, бо втішаєтесь ви, що спадщину Мою розграбовуєте, бо ви скачете, мов те теля по траві, та іржете, немов румаки...
JER|50|12|Збентежилася ваша мати занадто, застидалась родителька ваша... Оце для народів кінець: пустиня, сухоземля й степ!
JER|50|13|Від Господнього гніву вона незамешкана буде та стане спустошенням уся... Кожен, хто буде проходити повз Вавилон, остовпіє й засвище, як побачить усі ці порази його!
JER|50|14|Ушикуйтеся на Вавилон навкруги, всі, хто лука натягує! Стріляйте на нього, стріли не шкодуйте, бо він Господеві згрішив!
JER|50|15|Здійміть крик проти нього навколо! Він дав руку піддатись, стовпи його впали, зруйновані мури його, бо це помста Господня... Помстіться над ним: як зробив він зробіть так йому!
JER|50|16|Повигублюйте і сівача з Вавилону, і того, хто хапає серпа в часі жнив! Через меч переслідника вернуться всі до народу свого, і кожен до краю свого втече.
JER|50|17|Ізраїль вівця розпорошена, що леви погнали її: перший жер його цар асирійський, а останній цей Навуходоносор, цар вавилонський, розтрощив йому кості...
JER|50|18|Тому так промовляє Господь Саваот, Бог Ізраїлів: Ось Я покараю царя вавилонського й землю його, як Я покарав був царя асирійського.
JER|50|19|І верну Я Ізраїля на пасовисько його, і він пастися буде на Кармелі й Башані, і на горі на Єфремовій та на Ґілеаді душа його ситою буде.
JER|50|20|За тих днів й того часу говорить Господь будуть шукати провину Ізраїлеву, та не буде її, і прогріхи Юди, одначе не знайдені будуть вони, бо пробачу тому, кого Я позоставлю!
JER|50|21|На край Чварів подвійних, на нього піди й на мешканців Покарання! Поруйнуй і прокляттям вчини все за ними, говорить Господь, і зроби так усе, як тобі наказав!
JER|50|22|Гуркіт бою в краю та велике спустошення!
JER|50|23|Як побитий й поламаний молот всієї землі! Яким жахом зробивсь Вавилон для народів!
JER|50|24|Я пастку поставив на тебе, і схоплений ти, Вавилоне, хоча ти й не знав! Ти знайдений й схоплений був, бо ставав ти на прю проти Господа!
JER|50|25|Господь відчинив Своє сховище, і вийняв ізвідти знаряддя гніву Свого, це бо зайняття для Господа, Бога Саваота в халдейському краї.
JER|50|26|Ідіть ви на нього із краю землі, відчиніть його клуні, порозкладайте його, як снопи, і вчиніте закляттям його, хай не буде йому позосталого!
JER|50|27|Його всіх волів повбивайте, хай підуть вони на заріз! Горе їм, бо настав їхній день, час навіщення їх!
JER|50|28|Голос тих, що втікають і рятуються із вавилонського краю, щоб звістити на Сіоні про помсту Господа, нашого Бога, про помсту за храма Його.
JER|50|29|Скличте на Вавилона стрільців, усіх, хто лука натягує, табором станьте при ньому навколо, нехай йому втечі не буде! Відплатіте йому згідно з чином його, як зробив він зробіть так йому, бо гордим він став проти Господа, проти Святого Ізраїлевого!
JER|50|30|Тому то його юнаки всі поляжуть на площах його, а військові його того дня всі погинуть, говорить Господь.
JER|50|31|Ось Я проти тебе, о пихо, говорить Господь, Бог Саваот, бо день твій прийшов, час тебе покарати!
JER|50|32|І спіткнеться пиха й упаде, і не буде того, хто б підніс її. І огонь по містах його Я запалю, і він пожере всі довкілля його...
JER|50|33|Так говорить Господь Саваот: Сини Ізраїлеві й сини Юдині разом утискувані, і всі, що в полон їх забрали, тримають їх міцно, не хочуть їх випустити.
JER|50|34|Але Викупитель їх сильний, Господь Саваот Йому Ймення! Він конче розсудить їхню справу, щоб землю вспокоїти, а вавилонських мешканців стривожити.
JER|50|35|Меч на халдеїв, говорить Господь, і на мешканців Вавилону, і на князів його, і на його мудреців!
JER|50|36|Меч на ворожбитів і безглуздими стануть, меч на лицарство його і вони полякаються!
JER|50|37|Меч на коні його й на його колесниці, та на всю мішанину народів, яка серед нього, і стануть вони як жінки! Меч на скарби його й пограбовані будуть!
JER|50|38|Посуха на води його, й вони повисихають, бо це край божків, і шаліють вони від бовванів...
JER|50|39|Тому звірі пустинні там будуть сидіти з шакалами, і струсі будуть у ньому сидіти, і не буде заселений він вже навіки, і не буде замешканий він з роду в рід...
JER|50|40|Як Содом та Гоморру й сусідів її Бог був поруйнував, говорить Господь, так ніхто там не буде сидіти, і не буде в нім мешкати чужинцем син людський!
JER|50|41|Ось із півночі прийде народ, і люд великий, і численні царі, вони збуджені будуть із кінців землі:
JER|50|42|Лук та ратище міцно тримають, жорстокі вони й милосердя не мають, їхній голос, як море реве, вони їдуть на конях, на тебе вони вшикувались, як муж на війну, вавилонськая дочко!
JER|50|43|Почув цар вавилонський відомість про них, й опустилися руки йому, обхопив його страх і тремтіння, немов породіллю!...
JER|50|44|Ось підіймається він, немов лев, із темного лісу Йордану на водяні луки, і Я вмент зроблю, що він побіжить геть від них, а хто вибраний буде, того Я поставлю над ними! Бо хто є подібний Мені, і хто покличе Мене перед суд, і хто пастир такий, що перед обличчям Моїм він устоїть?
JER|50|45|Тому то послухайте задум Господній, що на Вавилон Він задумав, і думки Його ті, що на землю халдейську замислив: Поправді кажу вам, найменших з отари потягнуть, і попустошать пасовисько їхнє при них!
JER|50|46|Від розголосу про взяття Вавилону земля задрижить, і почується крик між народами!...
JER|51|1|Так говорить Господь: Ось Я бурю збуджу на отой Вавилон та на мешканців серця повстанців на Мене.
JER|51|2|І на Вавилон Я пошлю віяча, і розвіють його, і випорожнять його край, бо оточать його у день зла.
JER|51|3|Нехай лука свого напинає стрілець проти того, хто й собі напинає, проти того, хто своїм панцерем чваниться! І не змилуйтеся над його юнаками, закляттям учиніть усе військо його!
JER|51|4|І попадають вбиті в халдейському краї, і попробивані на його вулицях...
JER|51|5|Бо Ізраїль та Юда не вдівець він по Бозі своєму, по Господу Саваоту, та наповнився край їхній гріхом проти Святого Ізраїлевого.
JER|51|6|Утікайте з-серед Вавилону, і кожен урятовуйте душу свою! За провину його не погиньте, бо це Господеві час помсти, Він дасть відповідну заплату йому!
JER|51|7|Вавилон у Господній руці золотая це чаша, що всю землю напоювала: народи впивались вином тим його, тому пошаліли народи!
JER|51|8|Несподівано впав Вавилон і зруйнований він! Візьміте бальзаму для болю його, може буде загоєний він!
JER|51|9|Вавилон лікували, та він не був вилікуваний, покиньте його, і підемо кожен до краю свого, бо присуд його досягнув до небес, і дійшов аж до хмар!...
JER|51|10|Вивів Господь справедливості наші, прийдіть, і розповімо на Сіоні про чин оцей Господа, нашого Бога!
JER|51|11|Вигостріть стріли, візьміте щити! Збудив Господь духа мідійських царів, бо на Вавилон Його задум, понищити його, бо це помста Господня, помста за храма Його!
JER|51|12|Проти мурів Вавилону підійміте прапора, сторожу зміцніть, сторожів порозставляйте, і чати поставте, бо Господь і задумав, і зробив, що Він говорив був на мешканців Вавилону.
JER|51|13|О ти, що живеш над великими водами, що маєш скарбів багатенно, кінець твій прийшов, міра твоєї захланности!
JER|51|14|Господь Саваот присягав був душею Своєю: наповню людьми тебе, мов сараною, і на тебе вони крик військовий підіймуть!
JER|51|15|Своєю Він силою землю вчинив, Своєю премудрістю міцно поставив вселенну, і небо розтяг Своїм розумом.
JER|51|16|Як голос Його забринить, у небесах шумлять води, а коли підіймає Він хмари із краю землі, коли із дощем чинить блискавки та випроваджує вітер зо сховищ Своїх,
JER|51|17|тоді кожна людина в знанні туманіє, усяк золотар посоромлений через боввана, бо відлив його це неправда, і немає в них духа!
JER|51|18|Марнота вони, вони праця на сміх, в час навіщення їх вони згинуть!
JER|51|19|Не така, як оці, частка Яковова, бо все це Він створив, і Ізраїль племено спадщини Його, Господь Саваот Йому Ймення!
JER|51|20|Ти Мій молот, знаряддя військове, тобою поб'ю Я народи, і тобою Я вигублю царства!
JER|51|21|І тобою поб'ю Я коня й верхівця, і тобою поб'ю колесницю й її візника!
JER|51|22|І тобою поб'ю чоловіка та жінку, старого та хлопця тобою поб'ю, і тобою поб'ю юнака та дівчину!
JER|51|23|І тобою поб'ю пастуха й його стадо, і тобою поб'ю селянина та запряг його, і тобою поб'ю Я намісників та їхніх заступників!
JER|51|24|І Я відплачу Вавилонові і всім мешканцям халдеїв усе їхнє зло, що зробили в Сіоні на ваших очах, промовляє Господь!
JER|51|25|Оце Я на тебе, о горо ти згубна, говорить Господь, що всю землю ти губиш! І руку Свою простягну над тобою, і зо скель тебе скину, і зроблю горою горючою!
JER|51|26|І не братимуть з тебе наріжного каменя, ані каменя на підвалини, бо спустошенням вічним ти станеш, говорить Господь...
JER|51|27|Підійміте прапор на землі, засурміть у сурму між народами, приготуйте народи на бій проти нього, покличте на нього царства Арарату, Мінні та Ашкеназу, призначте гетьмана над ними, коней спровадьте, немов ту шорстку сарану!
JER|51|28|Приготуйте на бій проти нього народи, царів Мідії, намісників її та всіх її заступників, та ввесь край панування її!
JER|51|29|І затряслася земля, і корчитись стала від болю, бо здійснилися задуми Господа на Вавилон, щоб край вавилонський вчинити жахливим спустошенням та без мешканця...
JER|51|30|Силачі вавилонські воювати перестали, у твердинях осілись, загинула вся їхня сила, зробились, неначе жінки, оселі його попідпалювані, його засуви зламані...
JER|51|31|Бігун бігунові назустріч біжить, а посол назустріч послові, щоб звістити царю вавилонському, що з кінця до кінця взяте місто його,
JER|51|32|і броди захоплені, і фортеці огнем попалили, вояки перестрашені...
JER|51|33|Бо так промовляє Господь Саваот, Бог Ізраїлів: Дочка вавилонська мов тік в час топтання його: іще трохи й настане для неї час жнив!
JER|51|34|Пожер мене й стер мене Навуходоносор, цар вавилонський, поставив мене, як той посуд порожній, ковтнув він мене, немов змій, моїми розкошами сповнив свого живота, випхнув мене...
JER|51|35|Насилля моє й моє тіло на Вавилон, говорить мешканка Сіону, кров же моя на мешканців халдеїв, говорить Єрусалим!
JER|51|36|Тому так промовляє Господь: Оце Я змагаюсь за справу твою, і помщу твою помсту, і висушу море його, і джерело його висушу.
JER|51|37|І стане руїною цей Вавилон, мешканням шакалів, страхіттям та посміхом, і в ньому мешканця не буде!...
JER|51|38|Заревуть вони разом, немов левчуки, загарчать, немов ті левенята...
JER|51|39|Як вони порозпалюються, то зроблю їм бенкета та їх упою, щоб раділи й заснули сном вічним, і вже не пробудяться, каже Господь!
JER|51|40|Поспускаю Я їх, мов овець до зарізу, немов баранів із козлами.
JER|51|41|Як здобутий Шешах, і як схоплена слава всієї землі! Яким ось зробивсь Вавилон посеред народів!
JER|51|42|На Вавилон вийшло море, і вкрився він безліччю хвиль тих його.
JER|51|43|Міста його стануть спустошенням, краєм пустині та степу, тим краєм, що в ньому сидіти не буде ніяка людина, і не буде ходити по ньому син людський!
JER|51|44|І Я навіщу Бела в Вавилоні, і витягну з уст його те, що він був ковтнув, і вже народи до нього не будуть плисти, немов ріки, і мур вавилонський впаде!
JER|51|45|Мій народе, виходьте із нього й рятуйте від лютости гніву Господнього душу свою!
JER|51|46|І щоб серце ваше не слабло, а ви не злякалися вістки, почутої в краї, бо прийде цього року ця звістка, а потім того року та звістка, і буде насилля в краю, і повстане пануючий проти пануючого...
JER|51|47|Тому то ось дні настають, і навіщу Я божків Вавилону, і ввесь його край посоромлений буде, і всі його вбиті попадають в ньому!
JER|51|48|І над Вавилоном співатимуть небо й земля, і все, що є в них, бо на нього приходять спустошники з півночі, каже Господь.
JER|51|49|Вавилон мусить упасти за вбитих Ізраїлевих, як за Вавилон впали вбиті всієї землі...
JER|51|50|Хто втік від меча, ідіть, не ставайте! Пам'ятайте й здалека про Господа, а Єрусалим нехай буде на вашому серці!
JER|51|51|Застидалися ми, як почули цю ганьбу, сором покрив нам обличчя, бо чужинці прийшли у святиню Господнього дому...
JER|51|52|Тому то ось дні настають, говорить Господь, і бовванів його навіщу, і буде стогнати поранений по всім краї його!
JER|51|53|Коли б Вавилон аж до неба піднісся, і коли б уміцнив свою силу він на височині, то все таки прийдуть від Мене до нього спустошники, каже Господь!
JER|51|54|Чується крик з Вавилону, і велике понищення з краю халдеїв,
JER|51|55|бо пустошить Господь Вавилона і галас великий приглушує в ньому, і шумлять їхні хвилі, як води великі, і розлягається гуркіт їхнього голосу...
JER|51|56|Бо прийде спустошник на нього, на Вавилон, і схоплене буде лицарство його, їхній лук поламається, бож Бог відплати Господь, Він напевно заплатить!
JER|51|57|І впою його зверхників та мудреців його, намісників його та заступників його, і його лицарів, і сном вічним заснуть, і не збудяться, каже Цар, Господь Саваот Йому Ймення...
JER|51|58|Так говорить Господь Саваот: Товстий мур вавилонський аж до основ буде знищений, і брами високі його огнем будуть спалені, і мучились дармо народи, і для огню мордувались племена!...
JER|51|59|Слово, яке пророк Єремія наказав був Сераї, сину Нерійї, сина Махсеїного, коли він ішов з Седекією, Юдиним царем, до Вавилону, за четвертого року царювання його. А Серая був головним царським постельником.
JER|51|60|І написав Єремія все те лихо, що прийде на Вавилон, до однієї книги, усі ті слова, що написані на Вавилон.
JER|51|61|Я сказав Єремія до Сераї: Як прийдеш ти до Вавилону, то гляди, прочитай усі ці слова.
JER|51|62|І скажи: Господи, Ти провіщав на це місце, щоб вигубити його так, що не буде в ньому мешканця від людини й аж до скотини, бо буде воно спустошенням вічним.
JER|51|63|І станеться, як ти скінчиш читати цю книгу, прив'яжеш до неї каменя, і кинеш її до середини Ефрату,
JER|51|64|та й скажеш: Так потоне Вавилон, і не встане через те лихо, що Я на нього наведу, і вони попомучаться!... Аж досі слова Єремієні.
JER|52|1|Седекія був віку двадцяти й одного року, коли зацарював. А царював він в Єрусалимі одинадцять років; ім'я ж його матері Хамутал, дочка Єремії з Лівни.
JER|52|2|І робив він зло в Господніх очах, усе так, як робив був Єгояким.
JER|52|3|Бо через Господній гнів сталося це на Єрусалим та на Юду, аж поки Він не відкинув їх від Свого обличчя. А Седекія відпав від вавилонського царя.
JER|52|4|І сталося за дев'ятого року його царювання, десятого місяця, десятого дня місяця прийшов Навуходоносор, цар вавилонський, він та все військо його, на Єрусалим, і розтаборилися проти нього, і побудували проти нього вала навколо.
JER|52|5|І ввійшло місто в облогу аж до одинадцятого року царя Седекії.
JER|52|6|Четвертого місяця, дев'ятого дня місяця настав великий голод у місті, і не було хліба для народу краю.
JER|52|7|І пробитий був пролім у стіні міста, і всі вояки повтікали, і повиходили з міста вночі дорогою брами між двома мурами, що при царському садку, бо халдеї були при місті навколо. І пішли вони дорогою в степ.
JER|52|8|А халдейське військо погналося за царем, та й догнали Седекію в єрихонських степах, а все його військо розпорошилося від нього...
JER|52|9|І схопили царя, і відвели його до царя вавилонського до Рівли в краю Хамата, і там його той засудив.
JER|52|10|І цар вавилонський порізав Седекіїних синів на очах його, а також Юдиних зверхників він порізав у Рівлі...
JER|52|11|А очі Седекії він вибрав, і зв'язав його ланцюгами. І відвів його вавилонський цар до Вавилону, і посадив його до в'язниці аж до дня його смерти...
JER|52|12|А п'ятого місяця, десятого дня місяця, це дев'ятнадцятий рік царя Навуходоносора, вавилонського царя, прийшов до Єрусалиму Невузар'адан, начальник царської сторожі, що ставав перед обличчям вавилонського царя.
JER|52|13|І він спалив Господнього дома та дома царевого, і всі доми в Єрусалимі, і спалив кожного великого дома огнем.
JER|52|14|І мури навколо Єрусалиму порозбивало все халдейське військо, що було з начальником царської сторожі.
JER|52|15|А з бідноти народу та решту народу, що позостався в місті, і перебіжників, що перебігли до вавилонського царя, і решту простого люду повиганяв Невузар'адан, начальник царської сторожі.
JER|52|16|А з бідноти краю начальник царської сторожі позоставив декого за винарів та за рільників.
JER|52|17|А мідяні стовпи, що в Господньому домі, і підстави, і мідяне море, що в Господньому домі, халдеї поламали, і понесли всю їхню мідь до Вавилону.
JER|52|18|І горнята, і лопатки, і ножиці, і кропильниці, і ложки, і ввесь мідяний посуд, що ним служать, позабирали.
JER|52|19|І миски, і кадильниці, і кропильниці, і горнята, і свічники, і ложки, і жертовні миски, і що було золоте забрав золото, а що срібне срібло взяв начальник царської сторожі.
JER|52|20|Два стовпи, одне море, дванадцять мідяних волів, що під підставами, що цар Соломон поробив був для Господнього дому, не було й ваги для міді всіх цих речей!
JER|52|21|А стовпи вісімнадцять ліктів високість одного стовпа, і шнурок на дванадцять ліктів оточував його, а грубина його чотири пальці, всередині порожнявий.
JER|52|22|І маковиця на ньому мідяна, а високість однієї маковиці п'ять ліктів та мережка, і гранатові яблука на маковиці навколо, усе мідь. І для другого стовпа так само, і гранатові яблука.
JER|52|23|І було гранатових яблук дев'ятдесят і шість на кожну сторону, усіх гранатових яблук на мережці навколо сто.
JER|52|24|начальник царської сторожі взяв Сераю, головного священика, і Цефанію, другого священика, та трьох сторожів порога.
JER|52|25|А з міста взяв він одного евнуха, що був начальником над військовими, та семеро чоловіка з тих, що бачать цареве обличчя, що були знайдені в місті, і писаря, зверхника військового відділу, що записував народ краю до військового відділу, і шістдесят чоловіка з народу краю, що знаходилися в місті.
JER|52|26|І позабирав їх Невузар'адан, начальник царської сторожі, і відвів їх до вавилонського царя, до Рівли.
JER|52|27|І вдарив їх вавилонський цар, і позабивав їх у Рівлі, у хаматовому краї. І пішов Юда на вигнання з своєї землі!
JER|52|28|Оце той народ, що вигнав Навуходоносор: у сьомому році три тисячі й двадцять і три юдеї.
JER|52|29|У вісімнадцятому році Навуходоносора вигнав він з Єрусалиму вісім сотень тридцять і дві душі.
JER|52|30|У році двадцятому й третьому вигнав Невузар'адан, начальник царської сторожі, сім сотень сорок і п'ять душ юдеїв. Усіх душ чотири тисячі й шість сотень.
JER|52|31|І сталося за тридцятого й сьомого року вигнання Єгоякима, Юдиного царя, дванадцятого місяця, двадцятого й п'ятого дня місяця, Евіл-Меродах, цар вавилонський, у році свого зацарювання, змилувався над Єгоякимом, Юдиним царем, і вивів його з дому ув'язнення.
JER|52|32|І він говорив з ним добре, і поставив трона його понад трона царів, що були з ним у Вавилоні.
JER|52|33|І змінив в'язничну одежу його, і він завжди їв хліб перед ним по всі дні свого життя.
JER|52|34|А їжа його, їжа стала, видавалася йому від вавилонського царя, щоденне кожного дня, аж до дня його смерти, по всі дні його життя.
