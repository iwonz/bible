HAB|1|1|The oracle that Habakkuk the prophet saw.
HAB|1|2|O LORD, how long shall I cry for help, and you will not hear? Or cry to you "Violence!" and you will not save?
HAB|1|3|Why do you make me see iniquity, and why do you idly look at wrong? Destruction and violence are before me; strife and contention arise.
HAB|1|4|So the law is paralyzed, and justice never goes forth. For the wicked surround the righteous; so justice goes forth perverted.
HAB|1|5|"Look among the nations, and see; wonder and be astounded. For I am doing a work in your days that you would not believe if told.
HAB|1|6|For behold, I am raising up the Chaldeans, that bitter and hasty nation, who march through the breadth of the earth, to seize dwellings not their own.
HAB|1|7|They are dreaded and fearsome; their justice and dignity go forth from themselves.
HAB|1|8|Their horses are swifter than leopards, more fierce than the evening wolves; their horsemen press proudly on. Their horsemen come from afar; they fly like an eagle swift to devour.
HAB|1|9|They all come for violence, all their faces forward. They gather captives like sand.
HAB|1|10|At kings they scoff, and at rulers they laugh. They laugh at every fortress, for they pile up earth and take it.
HAB|1|11|Then they sweep by like the wind and go on, guilty men, whose own might is their god!"
HAB|1|12|Are you not from everlasting, O LORD my God, my Holy One? We shall not die. O LORD, you have ordained them as a judgment, and you, O Rock, have established them for reproof.
HAB|1|13|You who are of purer eyes than to see evil and cannot look at wrong, why do you idly look at traitors and are silent when the wicked swallows up the man more righteous than he?
HAB|1|14|You make mankind like the fish of the sea, like crawling things that have no ruler.
HAB|1|15|He brings all of them up with a hook; he drags them out with his net; he gathers them in his dragnet; so he rejoices and is glad.
HAB|1|16|Therefore he sacrifices to his net and makes offerings to his dragnet; for by them he lives in luxury, and his food is rich.
HAB|1|17|Is he then to keep on emptying his net and mercilessly killing nations forever?
HAB|2|1|I will take my stand at my watchpost and station myself on the tower, and look out to see what he will say to me, and what I will answer concerning my complaint.
HAB|2|2|And the LORD answered me: "Write the vision; make it plain on tablets, so he may run who reads it.
HAB|2|3|For still the vision awaits its appointed time; it hastens to the end- it will not lie. If it seems slow, wait for it; it will surely come; it will not delay.
HAB|2|4|"Behold, his soul is puffed up; it is not upright within him, but the righteous shall live by his faith.
HAB|2|5|"Moreover, wine is a traitor, an arrogant man who is never at rest. His greed is as wide as Sheol; like death he has never enough. He gathers for himself all nations and collects as his own all peoples."
HAB|2|6|Shall not all these take up their taunt against him, with scoffing and riddles for him, and say, "Woe to him who heaps up what is not his own- for how long?- and loads himself with pledges!"
HAB|2|7|Will not your debtors suddenly arise, and those awake who will make you tremble? Then you will be spoil for them.
HAB|2|8|Because you have plundered many nations, all the remnant of the peoples shall plunder you, for the blood of man and violence to the earth, to cities and all who dwell in them.
HAB|2|9|"Woe to him who gets evil gain for his house, to set his nest on high, to be safe from the reach of harm!
HAB|2|10|You have devised shame for your house by cutting off many peoples; you have forfeited your life.
HAB|2|11|For the stone will cry out from the wall, and the beam from the woodwork respond.
HAB|2|12|"Woe to him who builds a town with blood and founds a city on iniquity!
HAB|2|13|Behold, is it not from the LORD of hosts that peoples labor merely for fire, and nations weary themselves for nothing?
HAB|2|14|For the earth will be filled with the knowledge of the glory of the LORD as the waters cover the sea.
HAB|2|15|"Woe to him who makes his neighbors drink- you pour out your wrath and make them drunk, in order to gaze at their nakedness!
HAB|2|16|You will have your fill of shame instead of glory. Drink, yourself, and show your uncircumcision! The cup in the LORD'S right hand will come around to you, and utter shame will come upon your glory!
HAB|2|17|The violence done to Lebanon will overwhelm you, as will the destruction of the beasts that terrified them, for the blood of man and violence to the earth, to cities and all who dwell in them.
HAB|2|18|"What profit is an idol when its maker has shaped it, a metal image, a teacher of lies? For its maker trusts in his own creation when he makes speechless idols!
HAB|2|19|Woe to him who says to a wooden thing, Awake; to a silent stone, Arise! Can this teach? Behold, it is overlaid with gold and silver, and there is no breath at all in it.
HAB|2|20|But the LORD is in his holy temple; let all the earth keep silence before him."
HAB|3|1|A prayer of Habakkuk the prophet, according to Shigionoth.
HAB|3|2|O LORD, I have heard the report of you, and your work, O LORD, do I fear. In the midst of the years revive it; in the midst of the years make it known; in wrath remember mercy.
HAB|3|3|God came from Teman, and the Holy One from Mount Paran. His splendor covered the heavens, and the earth was full of his praise. Selah
HAB|3|4|His brightness was like the light; rays flashed from his hand; and there he veiled his power.
HAB|3|5|Before him went pestilence, and plague followed at his heels.
HAB|3|6|He stood and measured the earth; he looked and shook the nations; then the eternal mountains were scattered; the everlasting hills sank low. His were the everlasting ways.
HAB|3|7|I saw the tents of Cushan in affliction; the curtains of the land of Midian did tremble.
HAB|3|8|Was your wrath against the rivers, O LORD? Was your anger against the rivers, or your indignation against the sea, when you rode on your horses, on your chariot of salvation?
HAB|3|9|You stripped the sheath from your bow, calling for many arrows. Selah You split the earth with rivers.
HAB|3|10|The mountains saw you and writhed; the raging waters swept on; the deep gave forth its voice; it lifted its hands on high.
HAB|3|11|The sun and moon stood still in their place at the light of your arrows as they sped, at the flash of your glittering spear.
HAB|3|12|You marched through the earth in fury; you threshed the nations in anger.
HAB|3|13|You went out for the salvation of your people, for the salvation of your anointed. You crushed the head of the house of the wicked, laying him bare from thigh to neck. Selah
HAB|3|14|You pierced with his own arrows the heads of his warriors, who came like a whirlwind to scatter me, rejoicing as if to devour the poor in secret.
HAB|3|15|You trampled the sea with your horses, the surging of mighty waters.
HAB|3|16|I hear, and my body trembles; my lips quiver at the sound; rottenness enters into my bones; my legs tremble beneath me. Yet I will quietly wait for the day of trouble to come upon people who invade us.
HAB|3|17|Though the fig tree should not blossom, nor fruit be on the vines, the produce of the olive fail and the fields yield no food, the flock be cut off from the fold and there be no herd in the stalls,
HAB|3|18|yet I will rejoice in the LORD; I will take joy in the God of my salvation.
HAB|3|19|GOD, the Lord, is my strength; he makes my feet like the deer's; he makes me tread on my high places. To the choirmaster: with stringed instruments.
