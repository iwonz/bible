JUDG|1|1|Now after the death of Joshua it came to pass, that the children of Israel asked the LORD, saying, Who shall go up for us against the Canaanites first, to fight against them?
JUDG|1|2|And the LORD said, Judah shall go up: behold, I have delivered the land into his hand.
JUDG|1|3|And Judah said unto Simeon his brother, Come up with me into my lot, that we may fight against the Canaanites; and I likewise will go with thee into thy lot. So Simeon went with him.
JUDG|1|4|And Judah went up; and the LORD delivered the Canaanites and the Perizzites into their hand: and they slew of them in Bezek ten thousand men.
JUDG|1|5|And they found Adonibezek in Bezek: and they fought against him, and they slew the Canaanites and the Perizzites.
JUDG|1|6|But Adonibezek fled; and they pursued after him, and caught him, and cut off his thumbs and his great toes.
JUDG|1|7|And Adonibezek said, Threescore and ten kings, having their thumbs and their great toes cut off, gathered their meat under my table: as I have done, so God hath requited me. And they brought him to Jerusalem, and there he died.
JUDG|1|8|Now the children of Judah had fought against Jerusalem, and had taken it, and smitten it with the edge of the sword, and set the city on fire.
JUDG|1|9|And afterward the children of Judah went down to fight against the Canaanites, that dwelt in the mountain, and in the south, and in the valley.
JUDG|1|10|And Judah went against the Canaanites that dwelt in Hebron: (now the name of Hebron before was Kirjatharba:) and they slew Sheshai, and Ahiman, and Talmai.
JUDG|1|11|And from thence he went against the inhabitants of Debir: and the name of Debir before was Kirjathsepher:
JUDG|1|12|And Caleb said, He that smiteth Kirjathsepher, and taketh it, to him will I give Achsah my daughter to wife.
JUDG|1|13|And Othniel the son of Kenaz, Caleb's younger brother, took it: and he gave him Achsah his daughter to wife.
JUDG|1|14|And it came to pass, when she came to him, that she moved him to ask of her father a field: and she lighted from off her ass; and Caleb said unto her, What wilt thou?
JUDG|1|15|And she said unto him, Give me a blessing: for thou hast given me a south land; give me also springs of water. And Caleb gave her the upper springs and the nether springs.
JUDG|1|16|And the children of the Kenite, Moses' father in law, went up out of the city of palm trees with the children of Judah into the wilderness of Judah, which lieth in the south of Arad; and they went and dwelt among the people.
JUDG|1|17|And Judah went with Simeon his brother, and they slew the Canaanites that inhabited Zephath, and utterly destroyed it. And the name of the city was called Hormah.
JUDG|1|18|Also Judah took Gaza with the coast thereof, and Askelon with the coast thereof, and Ekron with the coast thereof.
JUDG|1|19|And the LORD was with Judah; and he drave out the inhabitants of the mountain; but could not drive out the inhabitants of the valley, because they had chariots of iron.
JUDG|1|20|And they gave Hebron unto Caleb, as Moses said: and he expelled thence the three sons of Anak.
JUDG|1|21|And the children of Benjamin did not drive out the Jebusites that inhabited Jerusalem; but the Jebusites dwell with the children of Benjamin in Jerusalem unto this day.
JUDG|1|22|And the house of Joseph, they also went up against Bethel: and the LORD was with them.
JUDG|1|23|And the house of Joseph sent to descry Bethel. (Now the name of the city before was Luz.)
JUDG|1|24|And the spies saw a man come forth out of the city, and they said unto him, Show us, we pray thee, the entrance into the city, and we will show thee mercy.
JUDG|1|25|And when he showed them the entrance into the city, they smote the city with the edge of the sword; but they let go the man and all his family.
JUDG|1|26|And the man went into the land of the Hittites, and built a city, and called the name thereof Luz: which is the name thereof unto this day.
JUDG|1|27|Neither did Manasseh drive out the inhabitants of Bethshean and her towns, nor Taanach and her towns, nor the inhabitants of Dor and her towns, nor the inhabitants of Ibleam and her towns, nor the inhabitants of Megiddo and her towns: but the Canaanites would dwell in that land.
JUDG|1|28|And it came to pass, when Israel was strong, that they put the Canaanites to tribute, and did not utterly drive them out.
JUDG|1|29|Neither did Ephraim drive out the Canaanites that dwelt in Gezer; but the Canaanites dwelt in Gezer among them.
JUDG|1|30|Neither did Zebulun drive out the inhabitants of Kitron, nor the inhabitants of Nahalol; but the Canaanites dwelt among them, and became tributaries.
JUDG|1|31|Neither did Asher drive out the inhabitants of Accho, nor the inhabitants of Zidon, nor of Ahlab, nor of Achzib, nor of Helbah, nor of Aphik, nor of Rehob:
JUDG|1|32|But the Asherites dwelt among the Canaanites, the inhabitants of the land: for they did not drive them out.
JUDG|1|33|Neither did Naphtali drive out the inhabitants of Bethshemesh, nor the inhabitants of Bethanath; but he dwelt among the Canaanites, the inhabitants of the land: nevertheless the inhabitants of Bethshemesh and of Bethanath became tributaries unto them.
JUDG|1|34|And the Amorites forced the children of Dan into the mountain: for they would not suffer them to come down to the valley:
JUDG|1|35|But the Amorites would dwell in mount Heres in Aijalon, and in Shaalbim: yet the hand of the house of Joseph prevailed, so that they became tributaries.
JUDG|1|36|And the coast of the Amorites was from the going up to Akrabbim, from the rock, and upward.
JUDG|2|1|And an angel of the LORD came up from Gilgal to Bochim, and said, I made you to go up out of Egypt, and have brought you unto the land which I sware unto your fathers; and I said, I will never break my covenant with you.
JUDG|2|2|And ye shall make no league with the inhabitants of this land; ye shall throw down their altars: but ye have not obeyed my voice: why have ye done this?
JUDG|2|3|Wherefore I also said, I will not drive them out from before you; but they shall be as thorns in your sides, and their gods shall be a snare unto you.
JUDG|2|4|And it came to pass, when the angel of the LORD spake these words unto all the children of Israel, that the people lifted up their voice, and wept.
JUDG|2|5|And they called the name of that place Bochim: and they sacrificed there unto the LORD.
JUDG|2|6|And when Joshua had let the people go, the children of Israel went every man unto his inheritance to possess the land.
JUDG|2|7|And the people served the LORD all the days of Joshua, and all the days of the elders that outlived Joshua, who had seen all the great works of the LORD, that he did for Israel.
JUDG|2|8|And Joshua the son of Nun, the servant of the LORD, died, being an hundred and ten years old.
JUDG|2|9|And they buried him in the border of his inheritance in Timnathheres, in the mount of Ephraim, on the north side of the hill Gaash.
JUDG|2|10|And also all that generation were gathered unto their fathers: and there arose another generation after them, which knew not the LORD, nor yet the works which he had done for Israel.
JUDG|2|11|And the children of Israel did evil in the sight of the LORD, and served Baalim:
JUDG|2|12|And they forsook the LORD God of their fathers, which brought them out of the land of Egypt, and followed other gods, of the gods of the people that were round about them, and bowed themselves unto them, and provoked the LORD to anger.
JUDG|2|13|And they forsook the LORD, and served Baal and Ashtaroth.
JUDG|2|14|And the anger of the LORD was hot against Israel, and he delivered them into the hands of spoilers that spoiled them, and he sold them into the hands of their enemies round about, so that they could not any longer stand before their enemies.
JUDG|2|15|Whithersoever they went out, the hand of the LORD was against them for evil, as the LORD had said, and as the LORD had sworn unto them: and they were greatly distressed.
JUDG|2|16|Nevertheless the LORD raised up judges, which delivered them out of the hand of those that spoiled them.
JUDG|2|17|And yet they would not hearken unto their judges, but they went a whoring after other gods, and bowed themselves unto them: they turned quickly out of the way which their fathers walked in, obeying the commandments of the LORD; but they did not so.
JUDG|2|18|And when the LORD raised them up judges, then the LORD was with the judge, and delivered them out of the hand of their enemies all the days of the judge: for it repented the LORD because of their groanings by reason of them that oppressed them and vexed them.
JUDG|2|19|And it came to pass, when the judge was dead, that they returned, and corrupted themselves more than their fathers, in following other gods to serve them, and to bow down unto them; they ceased not from their own doings, nor from their stubborn way.
JUDG|2|20|And the anger of the LORD was hot against Israel; and he said, Because that this people hath transgressed my covenant which I commanded their fathers, and have not hearkened unto my voice;
JUDG|2|21|I also will not henceforth drive out any from before them of the nations which Joshua left when he died:
JUDG|2|22|That through them I may prove Israel, whether they will keep the way of the LORD to walk therein, as their fathers did keep it, or not.
JUDG|2|23|Therefore the LORD left those nations, without driving them out hastily; neither delivered he them into the hand of Joshua.
JUDG|3|1|Now these are the nations which the LORD left, to prove Israel by them, even as many of Israel as had not known all the wars of Canaan;
JUDG|3|2|Only that the generations of the children of Israel might know, to teach them war, at the least such as before knew nothing thereof;
JUDG|3|3|Namely, five lords of the Philistines, and all the Canaanites, and the Sidonians, and the Hivites that dwelt in mount Lebanon, from mount Baalhermon unto the entering in of Hamath.
JUDG|3|4|And they were to prove Israel by them, to know whether they would hearken unto the commandments of the LORD, which he commanded their fathers by the hand of Moses.
JUDG|3|5|And the children of Israel dwelt among the Canaanites, Hittites, and Amorites, and Perizzites, and Hivites, and Jebusites:
JUDG|3|6|And they took their daughters to be their wives, and gave their daughters to their sons, and served their gods.
JUDG|3|7|And the children of Israel did evil in the sight of the LORD, and forgat the LORD their God, and served Baalim and the groves.
JUDG|3|8|Therefore the anger of the LORD was hot against Israel, and he sold them into the hand of Chushanrishathaim king of Mesopotamia: and the children of Israel served Chushanrishathaim eight years.
JUDG|3|9|And when the children of Israel cried unto the LORD, the LORD raised up a deliverer to the children of Israel, who delivered them, even Othniel the son of Kenaz, Caleb's younger brother.
JUDG|3|10|And the Spirit of the LORD came upon him, and he judged Israel, and went out to war: and the LORD delivered Chushanrishathaim king of Mesopotamia into his hand; and his hand prevailed against Chushanrishathaim.
JUDG|3|11|And the land had rest forty years. And Othniel the son of Kenaz died.
JUDG|3|12|And the children of Israel did evil again in the sight of the LORD: and the LORD strengthened Eglon the king of Moab against Israel, because they had done evil in the sight of the LORD.
JUDG|3|13|And he gathered unto him the children of Ammon and Amalek, and went and smote Israel, and possessed the city of palm trees.
JUDG|3|14|So the children of Israel served Eglon the king of Moab eighteen years.
JUDG|3|15|But when the children of Israel cried unto the LORD, the LORD raised them up a deliverer, Ehud the son of Gera, a Benjamite, a man lefthanded: and by him the children of Israel sent a present unto Eglon the king of Moab.
JUDG|3|16|But Ehud made him a dagger which had two edges, of a cubit length; and he did gird it under his raiment upon his right thigh.
JUDG|3|17|And he brought the present unto Eglon king of Moab: and Eglon was a very fat man.
JUDG|3|18|And when he had made an end to offer the present, he sent away the people that bare the present.
JUDG|3|19|But he himself turned again from the quarries that were by Gilgal, and said, I have a secret errand unto thee, O king: who said, Keep silence. And all that stood by him went out from him.
JUDG|3|20|And Ehud came unto him; and he was sitting in a summer parlor, which he had for himself alone. And Ehud said, I have a message from God unto thee. And he arose out of his seat.
JUDG|3|21|And Ehud put forth his left hand, and took the dagger from his right thigh, and thrust it into his belly:
JUDG|3|22|And the haft also went in after the blade; and the fat closed upon the blade, so that he could not draw the dagger out of his belly; and the dirt came out.
JUDG|3|23|Then Ehud went forth through the porch, and shut the doors of the parlor upon him, and locked them.
JUDG|3|24|When he was gone out, his servants came; and when they saw that, behold, the doors of the parlor were locked, they said, Surely he covereth his feet in his summer chamber.
JUDG|3|25|And they tarried till they were ashamed: and, behold, he opened not the doors of the parlor; therefore they took a key, and opened them: and, behold, their lord was fallen down dead on the earth.
JUDG|3|26|And Ehud escaped while they tarried, and passed beyond the quarries, and escaped unto Seirath.
JUDG|3|27|And it came to pass, when he was come, that he blew a trumpet in the mountain of Ephraim, and the children of Israel went down with him from the mount, and he before them.
JUDG|3|28|And he said unto them, Follow after me: for the LORD hath delivered your enemies the Moabites into your hand. And they went down after him, and took the fords of Jordan toward Moab, and suffered not a man to pass over.
JUDG|3|29|And they slew of Moab at that time about ten thousand men, all lusty, and all men of valor; and there escaped not a man.
JUDG|3|30|So Moab was subdued that day under the hand of Israel. And the land had rest fourscore years.
JUDG|3|31|And after him was Shamgar the son of Anath, which slew of the Philistines six hundred men with an ox goad: and he also delivered Israel.
JUDG|4|1|And the children of Israel again did evil in the sight of the LORD, when Ehud was dead.
JUDG|4|2|And the LORD sold them into the hand of Jabin king of Canaan, that reigned in Hazor; the captain of whose host was Sisera, which dwelt in Harosheth of the Gentiles.
JUDG|4|3|And the children of Israel cried unto the LORD: for he had nine hundred chariots of iron; and twenty years he mightily oppressed the children of Israel.
JUDG|4|4|And Deborah, a prophetess, the wife of Lapidoth, she judged Israel at that time.
JUDG|4|5|And she dwelt under the palm tree of Deborah between Ramah and Bethel in mount Ephraim: and the children of Israel came up to her for judgment.
JUDG|4|6|And she sent and called Barak the son of Abinoam out of Kedeshnaphtali, and said unto him, Hath not the LORD God of Israel commanded, saying, Go and draw toward mount Tabor, and take with thee ten thousand men of the children of Naphtali and of the children of Zebulun?
JUDG|4|7|And I will draw unto thee to the river Kishon Sisera, the captain of Jabin's army, with his chariots and his multitude; and I will deliver him into thine hand.
JUDG|4|8|And Barak said unto her, If thou wilt go with me, then I will go: but if thou wilt not go with me, then I will not go.
JUDG|4|9|And she said, I will surely go with thee: notwithstanding the journey that thou takest shall not be for thine honor; for the LORD shall sell Sisera into the hand of a woman. And Deborah arose, and went with Barak to Kedesh.
JUDG|4|10|And Barak called Zebulun and Naphtali to Kedesh; and he went up with ten thousand men at his feet: and Deborah went up with him.
JUDG|4|11|Now Heber the Kenite, which was of the children of Hobab the father in law of Moses, had severed himself from the Kenites, and pitched his tent unto the plain of Zaanaim, which is by Kedesh.
JUDG|4|12|And they showed Sisera that Barak the son of Abinoam was gone up to mount Tabor.
JUDG|4|13|And Sisera gathered together all his chariots, even nine hundred chariots of iron, and all the people that were with him, from Harosheth of the Gentiles unto the river of Kishon.
JUDG|4|14|And Deborah said unto Barak, Up; for this is the day in which the LORD hath delivered Sisera into thine hand: is not the LORD gone out before thee? So Barak went down from mount Tabor, and ten thousand men after him.
JUDG|4|15|And the LORD discomfited Sisera, and all his chariots, and all his host, with the edge of the sword before Barak; so that Sisera lighted down off his chariot, and fled away on his feet.
JUDG|4|16|But Barak pursued after the chariots, and after the host, unto Harosheth of the Gentiles: and all the host of Sisera fell upon the edge of the sword; and there was not a man left.
JUDG|4|17|Howbeit Sisera fled away on his feet to the tent of Jael the wife of Heber the Kenite: for there was peace between Jabin the king of Hazor and the house of Heber the Kenite.
JUDG|4|18|And Jael went out to meet Sisera, and said unto him, Turn in, my lord, turn in to me; fear not. And when he had turned in unto her into the tent, she covered him with a mantle.
JUDG|4|19|And he said unto her, Give me, I pray thee, a little water to drink; for I am thirsty. And she opened a bottle of milk, and gave him drink, and covered him.
JUDG|4|20|Again he said unto her, Stand in the door of the tent, and it shall be, when any man doth come and inquire of thee, and say, Is there any man here? that thou shalt say, No.
JUDG|4|21|Then Jael Heber's wife took a nail of the tent, and took an hammer in her hand, and went softly unto him, and smote the nail into his temples, and fastened it into the ground: for he was fast asleep and weary. So he died.
JUDG|4|22|And, behold, as Barak pursued Sisera, Jael came out to meet him, and said unto him, Come, and I will show thee the man whom thou seekest. And when he came into her tent, behold, Sisera lay dead, and the nail was in his temples.
JUDG|4|23|So God subdued on that day Jabin the king of Canaan before the children of Israel.
JUDG|4|24|And the hand of the children of Israel prospered, and prevailed against Jabin the king of Canaan, until they had destroyed Jabin king of Canaan.
JUDG|5|1|Then sang Deborah and Barak the son of Abinoam on that day, saying,
JUDG|5|2|Praise ye the LORD for the avenging of Israel, when the people willingly offered themselves.
JUDG|5|3|Hear, O ye kings; give ear, O ye princes; I, even I, will sing unto the LORD; I will sing praise to the LORD God of Israel.
JUDG|5|4|LORD, when thou wentest out of Seir, when thou marchedst out of the field of Edom, the earth trembled, and the heavens dropped, the clouds also dropped water.
JUDG|5|5|The mountains melted from before the LORD, even that Sinai from before the LORD God of Israel.
JUDG|5|6|In the days of Shamgar the son of Anath, in the days of Jael, the highways were unoccupied, and the travellers walked through byways.
JUDG|5|7|The inhabitants of the villages ceased, they ceased in Israel, until that I Deborah arose, that I arose a mother in Israel.
JUDG|5|8|They chose new gods; then was war in the gates: was there a shield or spear seen among forty thousand in Israel?
JUDG|5|9|My heart is toward the governors of Israel, that offered themselves willingly among the people. Bless ye the LORD.
JUDG|5|10|Speak, ye that ride on white asses, ye that sit in judgment, and walk by the way.
JUDG|5|11|They that are delivered from the noise of archers in the places of drawing water, there shall they rehearse the righteous acts of the LORD, even the righteous acts toward the inhabitants of his villages in Israel: then shall the people of the LORD go down to the gates.
JUDG|5|12|Awake, awake, Deborah: awake, awake, utter a song: arise, Barak, and lead thy captivity captive, thou son of Abinoam.
JUDG|5|13|Then he made him that remaineth have dominion over the nobles among the people: the LORD made me have dominion over the mighty.
JUDG|5|14|Out of Ephraim was there a root of them against Amalek; after thee, Benjamin, among thy people; out of Machir came down governors, and out of Zebulun they that handle the pen of the writer.
JUDG|5|15|And the princes of Issachar were with Deborah; even Issachar, and also Barak: he was sent on foot into the valley. For the divisions of Reuben there were great thoughts of heart.
JUDG|5|16|Why abodest thou among the sheepfolds, to hear the bleatings of the flocks? For the divisions of Reuben there were great searchings of heart.
JUDG|5|17|Gilead abode beyond Jordan: and why did Dan remain in ships? Asher continued on the sea shore, and abode in his breaches.
JUDG|5|18|Zebulun and Naphtali were a people that jeoparded their lives unto the death in the high places of the field.
JUDG|5|19|The kings came and fought, then fought the kings of Canaan in Taanach by the waters of Megiddo; they took no gain of money.
JUDG|5|20|They fought from heaven; the stars in their courses fought against Sisera.
JUDG|5|21|The river of Kishon swept them away, that ancient river, the river Kishon. O my soul, thou hast trodden down strength.
JUDG|5|22|Then were the horsehoofs broken by the means of the pransings, the pransings of their mighty ones.
JUDG|5|23|Curse ye Meroz, said the angel of the LORD, curse ye bitterly the inhabitants thereof; because they came not to the help of the LORD, to the help of the LORD against the mighty.
JUDG|5|24|Blessed above women shall Jael the wife of Heber the Kenite be, blessed shall she be above women in the tent.
JUDG|5|25|He asked water, and she gave him milk; she brought forth butter in a lordly dish.
JUDG|5|26|She put her hand to the nail, and her right hand to the workmen's hammer; and with the hammer she smote Sisera, she smote off his head, when she had pierced and stricken through his temples.
JUDG|5|27|At her feet he bowed, he fell, he lay down: at her feet he bowed, he fell: where he bowed, there he fell down dead.
JUDG|5|28|The mother of Sisera looked out at a window, and cried through the lattice, Why is his chariot so long in coming? why tarry the wheels of his chariots?
JUDG|5|29|Her wise ladies answered her, yea, she returned answer to herself,
JUDG|5|30|Have they not sped? have they not divided the prey; to every man a damsel or two; to Sisera a prey of divers colors, a prey of divers colors of needlework, of divers colors of needlework on both sides, meet for the necks of them that take the spoil?
JUDG|5|31|So let all thine enemies perish, O LORD: but let them that love him be as the sun when he goeth forth in his might. And the land had rest forty years.
JUDG|6|1|And the children of Israel did evil in the sight of the LORD: and the LORD delivered them into the hand of Midian seven years.
JUDG|6|2|And the hand of Midian prevailed against Israel: and because of the Midianites the children of Israel made them the dens which are in the mountains, and caves, and strong holds.
JUDG|6|3|And so it was, when Israel had sown, that the Midianites came up, and the Amalekites, and the children of the east, even they came up against them;
JUDG|6|4|And they encamped against them, and destroyed the increase of the earth, till thou come unto Gaza, and left no sustenance for Israel, neither sheep, nor ox, nor ass.
JUDG|6|5|For they came up with their cattle and their tents, and they came as grasshoppers for multitude; for both they and their camels were without number: and they entered into the land to destroy it.
JUDG|6|6|And Israel was greatly impoverished because of the Midianites; and the children of Israel cried unto the LORD.
JUDG|6|7|And it came to pass, when the children of Israel cried unto the LORD because of the Midianites,
JUDG|6|8|That the LORD sent a prophet unto the children of Israel, which said unto them, Thus saith the LORD God of Israel, I brought you up from Egypt, and brought you forth out of the house of bondage;
JUDG|6|9|And I delivered you out of the hand of the Egyptians, and out of the hand of all that oppressed you, and drave them out from before you, and gave you their land;
JUDG|6|10|And I said unto you, I am the LORD your God; fear not the gods of the Amorites, in whose land ye dwell: but ye have not obeyed my voice.
JUDG|6|11|And there came an angel of the LORD, and sat under an oak which was in Ophrah, that pertained unto Joash the Abiezrite: and his son Gideon threshed wheat by the winepress, to hide it from the Midianites.
JUDG|6|12|And the angel of the LORD appeared unto him, and said unto him, The LORD is with thee, thou mighty man of valor.
JUDG|6|13|And Gideon said unto him, Oh my Lord, if the LORD be with us, why then is all this befallen us? and where be all his miracles which our fathers told us of, saying, Did not the LORD bring us up from Egypt? but now the LORD hath forsaken us, and delivered us into the hands of the Midianites.
JUDG|6|14|And the LORD looked upon him, and said, Go in this thy might, and thou shalt save Israel from the hand of the Midianites: have not I sent thee?
JUDG|6|15|And he said unto him, Oh my Lord, wherewith shall I save Israel? behold, my family is poor in Manasseh, and I am the least in my father's house.
JUDG|6|16|And the LORD said unto him, Surely I will be with thee, and thou shalt smite the Midianites as one man.
JUDG|6|17|And he said unto him, If now I have found grace in thy sight, then show me a sign that thou talkest with me.
JUDG|6|18|Depart not hence, I pray thee, until I come unto thee, and bring forth my present, and set it before thee. And he said, I will tarry until thou come again.
JUDG|6|19|And Gideon went in, and made ready a kid, and unleavened cakes of an ephah of flour: the flesh he put in a basket, and he put the broth in a pot, and brought it out unto him under the oak, and presented it.
JUDG|6|20|And the angel of God said unto him, Take the flesh and the unleavened cakes, and lay them upon this rock, and pour out the broth. And he did so.
JUDG|6|21|Then the angel of the LORD put forth the end of the staff that was in his hand, and touched the flesh and the unleavened cakes; and there rose up fire out of the rock, and consumed the flesh and the unleavened cakes. Then the angel of the LORD departed out of his sight.
JUDG|6|22|And when Gideon perceived that he was an angel of the LORD, Gideon said, Alas, O LORD God! for because I have seen an angel of the LORD face to face.
JUDG|6|23|And the LORD said unto him, Peace be unto thee; fear not: thou shalt not die.
JUDG|6|24|Then Gideon built an altar there unto the LORD, and called it Jehovahshalom: unto this day it is yet in Ophrah of the Abiezrites.
JUDG|6|25|And it came to pass the same night, that the LORD said unto him, Take thy father's young bullock, even the second bullock of seven years old, and throw down the altar of Baal that thy father hath, and cut down the grove that is by it:
JUDG|6|26|And build an altar unto the LORD thy God upon the top of this rock, in the ordered place, and take the second bullock, and offer a burnt sacrifice with the wood of the grove which thou shalt cut down.
JUDG|6|27|Then Gideon took ten men of his servants, and did as the LORD had said unto him: and so it was, because he feared his father's household, and the men of the city, that he could not do it by day, that he did it by night.
JUDG|6|28|And when the men of the city arose early in the morning, behold, the altar of Baal was cast down, and the grove was cut down that was by it, and the second bullock was offered upon the altar that was built.
JUDG|6|29|And they said one to another, Who hath done this thing? And when they inquired and asked, they said, Gideon the son of Joash hath done this thing.
JUDG|6|30|Then the men of the city said unto Joash, Bring out thy son, that he may die: because he hath cast down the altar of Baal, and because he hath cut down the grove that was by it.
JUDG|6|31|And Joash said unto all that stood against him, Will ye plead for Baal? will ye save him? he that will plead for him, let him be put to death whilst it is yet morning: if he be a god, let him plead for himself, because one hath cast down his altar.
JUDG|6|32|Therefore on that day he called him Jerubbaal, saying, Let Baal plead against him, because he hath thrown down his altar.
JUDG|6|33|Then all the Midianites and the Amalekites and the children of the east were gathered together, and went over, and pitched in the valley of Jezreel.
JUDG|6|34|But the Spirit of the LORD came upon Gideon, and he blew a trumpet; and Abiezer was gathered after him.
JUDG|6|35|And he sent messengers throughout all Manasseh; who also was gathered after him: and he sent messengers unto Asher, and unto Zebulun, and unto Naphtali; and they came up to meet them.
JUDG|6|36|And Gideon said unto God, If thou wilt save Israel by mine hand, as thou hast said,
JUDG|6|37|Behold, I will put a fleece of wool in the floor; and if the dew be on the fleece only, and it be dry upon all the earth beside, then shall I know that thou wilt save Israel by mine hand, as thou hast said.
JUDG|6|38|And it was so: for he rose up early on the morrow, and thrust the fleece together, and wringed the dew out of the fleece, a bowl full of water.
JUDG|6|39|And Gideon said unto God, Let not thine anger be hot against me, and I will speak but this once: let me prove, I pray thee, but this once with the fleece; let it now be dry only upon the fleece, and upon all the ground let there be dew.
JUDG|6|40|And God did so that night: for it was dry upon the fleece only, and there was dew on all the ground.
JUDG|7|1|Then Jerubbaal, who is Gideon, and all the people that were with him, rose up early, and pitched beside the well of Harod: so that the host of the Midianites were on the north side of them, by the hill of Moreh, in the valley.
JUDG|7|2|And the LORD said unto Gideon, The people that are with thee are too many for me to give the Midianites into their hands, lest Israel vaunt themselves against me, saying, Mine own hand hath saved me.
JUDG|7|3|Now therefore go to, proclaim in the ears of the people, saying, Whosoever is fearful and afraid, let him return and depart early from mount Gilead. And there returned of the people twenty and two thousand; and there remained ten thousand.
JUDG|7|4|And the LORD said unto Gideon, The people are yet too many; bring them down unto the water, and I will try them for thee there: and it shall be, that of whom I say unto thee, This shall go with thee, the same shall go with thee; and of whomsoever I say unto thee, This shall not go with thee, the same shall not go.
JUDG|7|5|So he brought down the people unto the water: and the LORD said unto Gideon, Every one that lappeth of the water with his tongue, as a dog lappeth, him shalt thou set by himself; likewise every one that boweth down upon his knees to drink.
JUDG|7|6|And the number of them that lapped, putting their hand to their mouth, were three hundred men: but all the rest of the people bowed down upon their knees to drink water.
JUDG|7|7|And the LORD said unto Gideon, By the three hundred men that lapped will I save you, and deliver the Midianites into thine hand: and let all the other people go every man unto his place.
JUDG|7|8|So the people took victuals in their hand, and their trumpets: and he sent all the rest of Israel every man unto his tent, and retained those three hundred men: and the host of Midian was beneath him in the valley.
JUDG|7|9|And it came to pass the same night, that the LORD said unto him, Arise, get thee down unto the host; for I have delivered it into thine hand.
JUDG|7|10|But if thou fear to go down, go thou with Phurah thy servant down to the host:
JUDG|7|11|And thou shalt hear what they say; and afterward shall thine hands be strengthened to go down unto the host. Then went he down with Phurah his servant unto the outside of the armed men that were in the host.
JUDG|7|12|And the Midianites and the Amalekites and all the children of the east lay along in the valley like grasshoppers for multitude; and their camels were without number, as the sand by the sea side for multitude.
JUDG|7|13|And when Gideon was come, behold, there was a man that told a dream unto his fellow, and said, Behold, I dreamed a dream, and, lo, a cake of barley bread tumbled into the host of Midian, and came unto a tent, and smote it that it fell, and overturned it, that the tent lay along.
JUDG|7|14|And his fellow answered and said, This is nothing else save the sword of Gideon the son of Joash, a man of Israel: for into his hand hath God delivered Midian, and all the host.
JUDG|7|15|And it was so, when Gideon heard the telling of the dream, and the interpretation thereof, that he worshipped, and returned into the host of Israel, and said, Arise; for the LORD hath delivered into your hand the host of Midian.
JUDG|7|16|And he divided the three hundred men into three companies, and he put a trumpet in every man's hand, with empty pitchers, and lamps within the pitchers.
JUDG|7|17|And he said unto them, Look on me, and do likewise: and, behold, when I come to the outside of the camp, it shall be that, as I do, so shall ye do.
JUDG|7|18|When I blow with a trumpet, I and all that are with me, then blow ye the trumpets also on every side of all the camp, and say, The sword of the LORD, and of Gideon.
JUDG|7|19|So Gideon, and the hundred men that were with him, came unto the outside of the camp in the beginning of the middle watch; and they had but newly set the watch: and they blew the trumpets, and brake the pitchers that were in their hands.
JUDG|7|20|And the three companies blew the trumpets, and brake the pitchers, and held the lamps in their left hands, and the trumpets in their right hands to blow withal: and they cried, The sword of the LORD, and of Gideon.
JUDG|7|21|And they stood every man in his place round about the camp; and all the host ran, and cried, and fled.
JUDG|7|22|And the three hundred blew the trumpets, and the LORD set every man's sword against his fellow, even throughout all the host: and the host fled to Bethshittah in Zererath, and to the border of Abelmeholah, unto Tabbath.
JUDG|7|23|And the men of Israel gathered themselves together out of Naphtali, and out of Asher, and out of all Manasseh, and pursued after the Midianites.
JUDG|7|24|And Gideon sent messengers throughout all mount Ephraim, saying, come down against the Midianites, and take before them the waters unto Bethbarah and Jordan. Then all the men of Ephraim gathered themselves together, and took the waters unto Bethbarah and Jordan.
JUDG|7|25|And they took two princes of the Midianites, Oreb and Zeeb; and they slew Oreb upon the rock Oreb, and Zeeb they slew at the winepress of Zeeb, and pursued Midian, and brought the heads of Oreb and Zeeb to Gideon on the other side Jordan.
JUDG|8|1|And the men of Ephraim said unto him, Why hast thou served us thus, that thou calledst us not, when thou wentest to fight with the Midianites? And they did chide with him sharply.
JUDG|8|2|And he said unto them, What have I done now in comparison of you? Is not the gleaning of the grapes of Ephraim better than the vintage of Abiezer?
JUDG|8|3|God hath delivered into your hands the princes of Midian, Oreb and Zeeb: and what was I able to do in comparison of you? Then their anger was abated toward him, when he had said that.
JUDG|8|4|And Gideon came to Jordan, and passed over, he, and the three hundred men that were with him, faint, yet pursuing them.
JUDG|8|5|And he said unto the men of Succoth, Give, I pray you, loaves of bread unto the people that follow me; for they be faint, and I am pursuing after Zebah and Zalmunna, kings of Midian.
JUDG|8|6|And the princes of Succoth said, Are the hands of Zebah and Zalmunna now in thine hand, that we should give bread unto thine army?
JUDG|8|7|And Gideon said, Therefore when the LORD hath delivered Zebah and Zalmunna into mine hand, then I will tear your flesh with the thorns of the wilderness and with briers.
JUDG|8|8|And he went up thence to Penuel, and spake unto them likewise: and the men of Penuel answered him as the men of Succoth had answered him.
JUDG|8|9|And he spake also unto the men of Penuel, saying, When I come again in peace, I will break down this tower.
JUDG|8|10|Now Zebah and Zalmunna were in Karkor, and their hosts with them, about fifteen thousand men, all that were left of all the hosts of the children of the east: for there fell an hundred and twenty thousand men that drew sword.
JUDG|8|11|And Gideon went up by the way of them that dwelt in tents on the east of Nobah and Jogbehah, and smote the host; for the host was secure.
JUDG|8|12|And when Zebah and Zalmunna fled, he pursued after them, and took the two kings of Midian, Zebah and Zalmunna, and discomfited all the host.
JUDG|8|13|And Gideon the son of Joash returned from battle before the sun was up,
JUDG|8|14|And caught a young man of the men of Succoth, and inquired of him: and he described unto him the princes of Succoth, and the elders thereof, even threescore and seventeen men.
JUDG|8|15|And he came unto the men of Succoth, and said, Behold Zebah and Zalmunna, with whom ye did upbraid me, saying, Are the hands of Zebah and Zalmunna now in thine hand, that we should give bread unto thy men that are weary?
JUDG|8|16|And he took the elders of the city, and thorns of the wilderness and briers, and with them he taught the men of Succoth.
JUDG|8|17|And he beat down the tower of Penuel, and slew the men of the city.
JUDG|8|18|Then said he unto Zebah and Zalmunna, What manner of men were they whom ye slew at Tabor? And they answered, As thou art, so were they; each one resembled the children of a king.
JUDG|8|19|And he said, They were my brethren, even the sons of my mother: as the LORD liveth, if ye had saved them alive, I would not slay you.
JUDG|8|20|And he said unto Jether his firstborn, Up, and slay them. But the youth drew not his sword: for he feared, because he was yet a youth.
JUDG|8|21|Then Zebah and Zalmunna said, Rise thou, and fall upon us: for as the man is, so is his strength. And Gideon arose, and slew Zebah and Zalmunna, and took away the ornaments that were on their camels' necks.
JUDG|8|22|Then the men of Israel said unto Gideon, Rule thou over us, both thou, and thy son, and thy son's son also: for thou hast delivered us from the hand of Midian.
JUDG|8|23|And Gideon said unto them, I will not rule over you, neither shall my son rule over you: the LORD shall rule over you.
JUDG|8|24|And Gideon said unto them, I would desire a request of you, that ye would give me every man the earrings of his prey. (For they had golden earrings, because they were Ishmaelites.)
JUDG|8|25|And they answered, We will willingly give them. And they spread a garment, and did cast therein every man the earrings of his prey.
JUDG|8|26|And the weight of the golden earrings that he requested was a thousand and seven hundred shekels of gold; beside ornaments, and collars, and purple raiment that was on the kings of Midian, and beside the chains that were about their camels' necks.
JUDG|8|27|And Gideon made an ephod thereof, and put it in his city, even in Ophrah: and all Israel went thither a whoring after it: which thing became a snare unto Gideon, and to his house.
JUDG|8|28|Thus was Midian subdued before the children of Israel, so that they lifted up their heads no more. And the country was in quietness forty years in the days of Gideon.
JUDG|8|29|And Jerubbaal the son of Joash went and dwelt in his own house.
JUDG|8|30|And Gideon had threescore and ten sons of his body begotten: for he had many wives.
JUDG|8|31|And his concubine that was in Shechem, she also bare him a son, whose name he called Abimelech.
JUDG|8|32|And Gideon the son of Joash died in a good old age, and was buried in the sepulchre of Joash his father, in Ophrah of the Abiezrites.
JUDG|8|33|And it came to pass, as soon as Gideon was dead, that the children of Israel turned again, and went a whoring after Baalim, and made Baalberith their god.
JUDG|8|34|And the children of Israel remembered not the LORD their God, who had delivered them out of the hands of all their enemies on every side:
JUDG|8|35|Neither showed they kindness to the house of Jerubbaal, namely, Gideon, according to all the goodness which he had showed unto Israel.
JUDG|9|1|And Abimelech the son of Jerubbaal went to Shechem unto his mother's brethren, and communed with them, and with all the family of the house of his mother's father, saying,
JUDG|9|2|Speak, I pray you, in the ears of all the men of Shechem, Whether is better for you, either that all the sons of Jerubbaal, which are threescore and ten persons, reign over you, or that one reign over you? remember also that I am your bone and your flesh.
JUDG|9|3|And his mother's brethren spake of him in the ears of all the men of Shechem all these words: and their hearts inclined to follow Abimelech; for they said, He is our brother.
JUDG|9|4|And they gave him threescore and ten pieces of silver out of the house of Baalberith, wherewith Abimelech hired vain and light persons, which followed him.
JUDG|9|5|And he went unto his father's house at Ophrah, and slew his brethren the sons of Jerubbaal, being threescore and ten persons, upon one stone: notwithstanding yet Jotham the youngest son of Jerubbaal was left; for he hid himself.
JUDG|9|6|And all the men of Shechem gathered together, and all the house of Millo, and went, and made Abimelech king, by the plain of the pillar that was in Shechem.
JUDG|9|7|And when they told it to Jotham, he went and stood in the top of mount Gerizim, and lifted up his voice, and cried, and said unto them, Hearken unto me, ye men of Shechem, that God may hearken unto you.
JUDG|9|8|The trees went forth on a time to anoint a king over them; and they said unto the olive tree, Reign thou over us.
JUDG|9|9|But the olive tree said unto them, Should I leave my fatness, wherewith by me they honor God and man, and go to be promoted over the trees?
JUDG|9|10|And the trees said to the fig tree, Come thou, and reign over us.
JUDG|9|11|But the fig tree said unto them, Should I forsake my sweetness, and my good fruit, and go to be promoted over the trees?
JUDG|9|12|Then said the trees unto the vine, Come thou, and reign over us.
JUDG|9|13|And the vine said unto them, Should I leave my wine, which cheereth God and man, and go to be promoted over the trees?
JUDG|9|14|Then said all the trees unto the bramble, Come thou, and reign over us.
JUDG|9|15|And the bramble said unto the trees, If in truth ye anoint me king over you, then come and put your trust in my shadow: and if not, let fire come out of the bramble, and devour the cedars of Lebanon.
JUDG|9|16|Now therefore, if ye have done truly and sincerely, in that ye have made Abimelech king, and if ye have dealt well with Jerubbaal and his house, and have done unto him according to the deserving of his hands;
JUDG|9|17|(For my father fought for you, and adventured his life far, and delivered you out of the hand of Midian:
JUDG|9|18|And ye are risen up against my father's house this day, and have slain his sons, threescore and ten persons, upon one stone, and have made Abimelech, the son of his maidservant, king over the men of Shechem, because he is your brother;)
JUDG|9|19|If ye then have dealt truly and sincerely with Jerubbaal and with his house this day, then rejoice ye in Abimelech, and let him also rejoice in you:
JUDG|9|20|But if not, let fire come out from Abimelech, and devour the men of Shechem, and the house of Millo; and let fire come out from the men of Shechem, and from the house of Millo, and devour Abimelech.
JUDG|9|21|And Jotham ran away, and fled, and went to Beer, and dwelt there, for fear of Abimelech his brother.
JUDG|9|22|When Abimelech had reigned three years over Israel,
JUDG|9|23|Then God sent an evil spirit between Abimelech and the men of Shechem; and the men of Shechem dealt treacherously with Abimelech:
JUDG|9|24|That the cruelty done to the threescore and ten sons of Jerubbaal might come, and their blood be laid upon Abimelech their brother, which slew them; and upon the men of Shechem, which aided him in the killing of his brethren.
JUDG|9|25|And the men of Shechem set liers in wait for him in the top of the mountains, and they robbed all that came along that way by them: and it was told Abimelech.
JUDG|9|26|And Gaal the son of Ebed came with his brethren, and went over to Shechem: and the men of Shechem put their confidence in him.
JUDG|9|27|And they went out into the fields, and gathered their vineyards, and trode the grapes, and made merry, and went into the house of their god, and did eat and drink, and cursed Abimelech.
JUDG|9|28|And Gaal the son of Ebed said, Who is Abimelech, and who is Shechem, that we should serve him? is not he the son of Jerubbaal? and Zebul his officer? serve the men of Hamor the father of Shechem: for why should we serve him?
JUDG|9|29|And would to God this people were under my hand! then would I remove Abimelech. And he said to Abimelech, Increase thine army, and come out.
JUDG|9|30|And when Zebul the ruler of the city heard the words of Gaal the son of Ebed, his anger was kindled.
JUDG|9|31|And he sent messengers unto Abimelech privily, saying, Behold, Gaal the son of Ebed and his brethren be come to Shechem; and, behold, they fortify the city against thee.
JUDG|9|32|Now therefore up by night, thou and the people that is with thee, and lie in wait in the field:
JUDG|9|33|And it shall be, that in the morning, as soon as the sun is up, thou shalt rise early, and set upon the city: and, behold, when he and the people that is with him come out against thee, then mayest thou do to them as thou shalt find occasion.
JUDG|9|34|And Abimelech rose up, and all the people that were with him, by night, and they laid wait against Shechem in four companies.
JUDG|9|35|And Gaal the son of Ebed went out, and stood in the entering of the gate of the city: and Abimelech rose up, and the people that were with him, from lying in wait.
JUDG|9|36|And when Gaal saw the people, he said to Zebul, Behold, there come people down from the top of the mountains. And Zebul said unto him, Thou seest the shadow of the mountains as if they were men.
JUDG|9|37|And Gaal spake again, and said, See there come people down by the middle of the land, and another company come along by the plain of Meonenim.
JUDG|9|38|Then said Zebul unto him, Where is now thy mouth, wherewith thou saidst, Who is Abimelech, that we should serve him? is not this the people that thou hast despised? go out, I pray now, and fight with them.
JUDG|9|39|And Gaal went out before the men of Shechem, and fought with Abimelech.
JUDG|9|40|And Abimelech chased him, and he fled before him, and many were overthrown and wounded, even unto the entering of the gate.
JUDG|9|41|And Abimelech dwelt at Arumah: and Zebul thrust out Gaal and his brethren, that they should not dwell in Shechem.
JUDG|9|42|And it came to pass on the morrow, that the people went out into the field; and they told Abimelech.
JUDG|9|43|And he took the people, and divided them into three companies, and laid wait in the field, and looked, and, behold, the people were come forth out of the city; and he rose up against them, and smote them.
JUDG|9|44|And Abimelech, and the company that was with him, rushed forward, and stood in the entering of the gate of the city: and the two other companies ran upon all the people that were in the fields, and slew them.
JUDG|9|45|And Abimelech fought against the city all that day; and he took the city, and slew the people that was therein, and beat down the city, and sowed it with salt.
JUDG|9|46|And when all the men of the tower of Shechem heard that, they entered into an hold of the house of the god Berith.
JUDG|9|47|And it was told Abimelech, that all the men of the tower of Shechem were gathered together.
JUDG|9|48|And Abimelech gat him up to mount Zalmon, he and all the people that were with him; and Abimelech took an axe in his hand, and cut down a bough from the trees, and took it, and laid it on his shoulder, and said unto the people that were with him, What ye have seen me do, make haste, and do as I have done.
JUDG|9|49|And all the people likewise cut down every man his bough, and followed Abimelech, and put them to the hold, and set the hold on fire upon them; so that all the men of the tower of Shechem died also, about a thousand men and women.
JUDG|9|50|Then went Abimelech to Thebez, and encamped against Thebez, and took it.
JUDG|9|51|But there was a strong tower within the city, and thither fled all the men and women, and all they of the city, and shut it to them, and gat them up to the top of the tower.
JUDG|9|52|And Abimelech came unto the tower, and fought against it, and went hard unto the door of the tower to burn it with fire.
JUDG|9|53|And a certain woman cast a piece of a millstone upon Abimelech's head, and all to brake his skull.
JUDG|9|54|Then he called hastily unto the young man his armourbearer, and said unto him, Draw thy sword, and slay me, that men say not of me, A women slew him. And his young man thrust him through, and he died.
JUDG|9|55|And when the men of Israel saw that Abimelech was dead, they departed every man unto his place.
JUDG|9|56|Thus God rendered the wickedness of Abimelech, which he did unto his father, in slaying his seventy brethren:
JUDG|9|57|And all the evil of the men of Shechem did God render upon their heads: and upon them came the curse of Jotham the son of Jerubbaal.
JUDG|10|1|And after Abimelech there arose to defend Israel Tola the son of Puah, the son of Dodo, a man of Issachar; and he dwelt in Shamir in mount Ephraim.
JUDG|10|2|And he judged Israel twenty and three years, and died, and was buried in Shamir.
JUDG|10|3|And after him arose Jair, a Gileadite, and judged Israel twenty and two years.
JUDG|10|4|And he had thirty sons that rode on thirty ass colts, and they had thirty cities, which are called Havothjair unto this day, which are in the land of Gilead.
JUDG|10|5|And Jair died, and was buried in Camon.
JUDG|10|6|And the children of Israel did evil again in the sight of the LORD, and served Baalim, and Ashtaroth, and the gods of Syria, and the gods of Zidon, and the gods of Moab, and the gods of the children of Ammon, and the gods of the Philistines, and forsook the LORD, and served not him.
JUDG|10|7|And the anger of the LORD was hot against Israel, and he sold them into the hands of the Philistines, and into the hands of the children of Ammon.
JUDG|10|8|And that year they vexed and oppressed the children of Israel: eighteen years, all the children of Israel that were on the other side Jordan in the land of the Amorites, which is in Gilead.
JUDG|10|9|Moreover the children of Ammon passed over Jordan to fight also against Judah, and against Benjamin, and against the house of Ephraim; so that Israel was sore distressed.
JUDG|10|10|And the children of Israel cried unto the LORD, saying, We have sinned against thee, both because we have forsaken our God, and also served Baalim.
JUDG|10|11|And the LORD said unto the children of Israel, Did not I deliver you from the Egyptians, and from the Amorites, from the children of Ammon, and from the Philistines?
JUDG|10|12|The Zidonians also, and the Amalekites, and the Maonites, did oppress you; and ye cried to me, and I delivered you out of their hand.
JUDG|10|13|Yet ye have forsaken me, and served other gods: wherefore I will deliver you no more.
JUDG|10|14|Go and cry unto the gods which ye have chosen; let them deliver you in the time of your tribulation.
JUDG|10|15|And the children of Israel said unto the LORD, We have sinned: do thou unto us whatsoever seemeth good unto thee; deliver us only, we pray thee, this day.
JUDG|10|16|And they put away the strange gods from among them, and served the LORD: and his soul was grieved for the misery of Israel.
JUDG|10|17|Then the children of Ammon were gathered together, and encamped in Gilead. And the children of Israel assembled themselves together, and encamped in Mizpeh.
JUDG|10|18|And the people and princes of Gilead said one to another, What man is he that will begin to fight against the children of Ammon? he shall be head over all the inhabitants of Gilead.
JUDG|11|1|Now Jephthah the Gileadite was a mighty man of valor, and he was the son of an harlot: and Gilead begat Jephthah.
JUDG|11|2|And Gilead's wife bare him sons; and his wife's sons grew up, and they thrust out Jephthah, and said unto him, Thou shalt not inherit in our father's house; for thou art the son of a strange woman.
JUDG|11|3|Then Jephthah fled from his brethren, and dwelt in the land of Tob: and there were gathered vain men to Jephthah, and went out with him.
JUDG|11|4|And it came to pass in process of time, that the children of Ammon made war against Israel.
JUDG|11|5|And it was so, that when the children of Ammon made war against Israel, the elders of Gilead went to fetch Jephthah out of the land of Tob:
JUDG|11|6|And they said unto Jephthah, Come, and be our captain, that we may fight with the children of Ammon.
JUDG|11|7|And Jephthah said unto the elders of Gilead, Did not ye hate me, and expel me out of my father's house? and why are ye come unto me now when ye are in distress?
JUDG|11|8|And the elders of Gilead said unto Jephthah, Therefore we turn again to thee now, that thou mayest go with us, and fight against the children of Ammon, and be our head over all the inhabitants of Gilead.
JUDG|11|9|And Jephthah said unto the elders of Gilead, If ye bring me home again to fight against the children of Ammon, and the LORD deliver them before me, shall I be your head?
JUDG|11|10|And the elders of Gilead said unto Jephthah, The LORD be witness between us, if we do not so according to thy words.
JUDG|11|11|Then Jephthah went with the elders of Gilead, and the people made him head and captain over them: and Jephthah uttered all his words before the LORD in Mizpeh.
JUDG|11|12|And Jephthah sent messengers unto the king of the children of Ammon, saying, What hast thou to do with me, that thou art come against me to fight in my land?
JUDG|11|13|And the king of the children of Ammon answered unto the messengers of Jephthah, Because Israel took away my land, when they came up out of Egypt, from Arnon even unto Jabbok, and unto Jordan: now therefore restore those lands again peaceably.
JUDG|11|14|And Jephthah sent messengers again unto the king of the children of Ammon:
JUDG|11|15|And said unto him, Thus saith Jephthah, Israel took not away the land of Moab, nor the land of the children of Ammon:
JUDG|11|16|But when Israel came up from Egypt, and walked through the wilderness unto the Red sea, and came to Kadesh;
JUDG|11|17|Then Israel sent messengers unto the king of Edom, saying, Let me, I pray thee, pass through thy land: but the king of Edom would not hearken thereto. And in like manner they sent unto the king of Moab: but he would not consent: and Israel abode in Kadesh.
JUDG|11|18|Then they went along through the wilderness, and compassed the land of Edom, and the land of Moab, and came by the east side of the land of Moab, and pitched on the other side of Arnon, but came not within the border of Moab: for Arnon was the border of Moab.
JUDG|11|19|And Israel sent messengers unto Sihon king of the Amorites, the king of Heshbon; and Israel said unto him, Let us pass, we pray thee, through thy land into my place.
JUDG|11|20|But Sihon trusted not Israel to pass through his coast: but Sihon gathered all his people together, and pitched in Jahaz, and fought against Israel.
JUDG|11|21|And the LORD God of Israel delivered Sihon and all his people into the hand of Israel, and they smote them: so Israel possessed all the land of the Amorites, the inhabitants of that country.
JUDG|11|22|And they possessed all the coasts of the Amorites, from Arnon even unto Jabbok, and from the wilderness even unto Jordan.
JUDG|11|23|So now the LORD God of Israel hath dispossessed the Amorites from before his people Israel, and shouldest thou possess it?
JUDG|11|24|Wilt not thou possess that which Chemosh thy god giveth thee to possess? So whomsoever the LORD our God shall drive out from before us, them will we possess.
JUDG|11|25|And now art thou any thing better than Balak the son of Zippor, king of Moab? did he ever strive against Israel, or did he ever fight against them,
JUDG|11|26|While Israel dwelt in Heshbon and her towns, and in Aroer and her towns, and in all the cities that be along by the coasts of Arnon, three hundred years? why therefore did ye not recover them within that time?
JUDG|11|27|Wherefore I have not sinned against thee, but thou doest me wrong to war against me: the LORD the Judge be judge this day between the children of Israel and the children of Ammon.
JUDG|11|28|Howbeit the king of the children of Ammon hearkened not unto the words of Jephthah which he sent him.
JUDG|11|29|Then the Spirit of the LORD came upon Jephthah, and he passed over Gilead, and Manasseh, and passed over Mizpeh of Gilead, and from Mizpeh of Gilead he passed over unto the children of Ammon.
JUDG|11|30|And Jephthah vowed a vow unto the LORD, and said, If thou shalt without fail deliver the children of Ammon into mine hands,
JUDG|11|31|Then it shall be, that whatsoever cometh forth of the doors of my house to meet me, when I return in peace from the children of Ammon, shall surely be the LORD's, and I will offer it up for a burnt offering.
JUDG|11|32|So Jephthah passed over unto the children of Ammon to fight against them; and the LORD delivered them into his hands.
JUDG|11|33|And he smote them from Aroer, even till thou come to Minnith, even twenty cities, and unto the plain of the vineyards, with a very great slaughter. Thus the children of Ammon were subdued before the children of Israel.
JUDG|11|34|And Jephthah came to Mizpeh unto his house, and, behold, his daughter came out to meet him with timbrels and with dances: and she was his only child; beside her he had neither son nor daughter.
JUDG|11|35|And it came to pass, when he saw her, that he rent his clothes, and said, Alas, my daughter! thou hast brought me very low, and thou art one of them that trouble me: for I have opened my mouth unto the LORD, and I cannot go back.
JUDG|11|36|And she said unto him, My father, if thou hast opened thy mouth unto the LORD, do to me according to that which hath proceeded out of thy mouth; forasmuch as the LORD hath taken vengeance for thee of thine enemies, even of the children of Ammon.
JUDG|11|37|And she said unto her father, Let this thing be done for me: let me alone two months, that I may go up and down upon the mountains, and bewail my virginity, I and my fellows.
JUDG|11|38|And he said, Go. And he sent her away for two months: and she went with her companions, and bewailed her virginity upon the mountains.
JUDG|11|39|And it came to pass at the end of two months, that she returned unto her father, who did with her according to his vow which he had vowed: and she knew no man. And it was a custom in Israel,
JUDG|11|40|That the daughters of Israel went yearly to lament the daughter of Jephthah the Gileadite four days in a year.
JUDG|12|1|And the men of Ephraim gathered themselves together, and went northward, and said unto Jephthah, Wherefore passedst thou over to fight against the children of Ammon, and didst not call us to go with thee? we will burn thine house upon thee with fire.
JUDG|12|2|And Jephthah said unto them, I and my people were at great strife with the children of Ammon; and when I called you, ye delivered me not out of their hands.
JUDG|12|3|And when I saw that ye delivered me not, I put my life in my hands, and passed over against the children of Ammon, and the LORD delivered them into my hand: wherefore then are ye come up unto me this day, to fight against me?
JUDG|12|4|Then Jephthah gathered together all the men of Gilead, and fought with Ephraim: and the men of Gilead smote Ephraim, because they said, Ye Gileadites are fugitives of Ephraim among the Ephraimites, and among the Manassites.
JUDG|12|5|And the Gileadites took the passages of Jordan before the Ephraimites: and it was so, that when those Ephraimites which were escaped said, Let me go over; that the men of Gilead said unto him, Art thou an Ephraimite? If he said, Nay;
JUDG|12|6|Then said they unto him, Say now Shibboleth: and he said Sibboleth: for he could not frame to pronounce it right. Then they took him, and slew him at the passages of Jordan: and there fell at that time of the Ephraimites forty and two thousand.
JUDG|12|7|And Jephthah judged Israel six years. Then died Jephthah the Gileadite, and was buried in one of the cities of Gilead.
JUDG|12|8|And after him Ibzan of Bethlehem judged Israel.
JUDG|12|9|And he had thirty sons, and thirty daughters, whom he sent abroad, and took in thirty daughters from abroad for his sons. And he judged Israel seven years.
JUDG|12|10|Then died Ibzan, and was buried at Bethlehem.
JUDG|12|11|And after him Elon, a Zebulonite, judged Israel; and he judged Israel ten years.
JUDG|12|12|And Elon the Zebulonite died, and was buried in Aijalon in the country of Zebulun.
JUDG|12|13|And after him Abdon the son of Hillel, a Pirathonite, judged Israel.
JUDG|12|14|And he had forty sons and thirty nephews, that rode on threescore and ten ass colts: and he judged Israel eight years.
JUDG|12|15|And Abdon the son of Hillel the Pirathonite died, and was buried in Pirathon in the land of Ephraim, in the mount of the Amalekites.
JUDG|13|1|And the children of Israel did evil again in the sight of the LORD; and the LORD delivered them into the hand of the Philistines forty years.
JUDG|13|2|And there was a certain man of Zorah, of the family of the Danites, whose name was Manoah; and his wife was barren, and bare not.
JUDG|13|3|And the angel of the LORD appeared unto the woman, and said unto her, Behold now, thou art barren, and bearest not: but thou shalt conceive, and bear a son.
JUDG|13|4|Now therefore beware, I pray thee, and drink not wine nor strong drink, and eat not any unclean thing:
JUDG|13|5|For, lo, thou shalt conceive, and bear a son; and no razor shall come on his head: for the child shall be a Nazarite unto God from the womb: and he shall begin to deliver Israel out of the hand of the Philistines.
JUDG|13|6|Then the woman came and told her husband, saying, A man of God came unto me, and his countenance was like the countenance of an angel of God, very terrible: but I asked him not whence he was, neither told he me his name:
JUDG|13|7|But he said unto me, Behold, thou shalt conceive, and bear a son; and now drink no wine nor strong drink, neither eat any unclean thing: for the child shall be a Nazarite to God from the womb to the day of his death.
JUDG|13|8|Then Manoah intreated the LORD, and said, O my Lord, let the man of God which thou didst send come again unto us, and teach us what we shall do unto the child that shall be born.
JUDG|13|9|And God hearkened to the voice of Manoah; and the angel of God came again unto the woman as she sat in the field: but Manoah her husband was not with her.
JUDG|13|10|And the woman made haste, and ran, and showed her husband, and said unto him, Behold, the man hath appeared unto me, that came unto me the other day.
JUDG|13|11|And Manoah arose, and went after his wife, and came to the man, and said unto him, Art thou the man that spakest unto the woman? And he said, I am.
JUDG|13|12|And Manoah said, Now let thy words come to pass. How shall we order the child, and how shall we do unto him?
JUDG|13|13|And the angel of the LORD said unto Manoah, Of all that I said unto the woman let her beware.
JUDG|13|14|She may not eat of any thing that cometh of the vine, neither let her drink wine or strong drink, nor eat any unclean thing: all that I commanded her let her observe.
JUDG|13|15|And Manoah said unto the angel of the LORD, I pray thee, let us detain thee, until we shall have made ready a kid for thee.
JUDG|13|16|And the angel of the LORD said unto Manoah, Though thou detain me, I will not eat of thy bread: and if thou wilt offer a burnt offering, thou must offer it unto the LORD. For Manoah knew not that he was an angel of the LORD.
JUDG|13|17|And Manoah said unto the angel of the LORD, What is thy name, that when thy sayings come to pass we may do thee honor?
JUDG|13|18|And the angel of the LORD said unto him, Why askest thou thus after my name, seeing it is secret?
JUDG|13|19|So Manoah took a kid with a meat offering, and offered it upon a rock unto the LORD: and the angel did wonderously; and Manoah and his wife looked on.
JUDG|13|20|For it came to pass, when the flame went up toward heaven from off the altar, that the angel of the LORD ascended in the flame of the altar. And Manoah and his wife looked on it, and fell on their faces to the ground.
JUDG|13|21|But the angel of the LORD did no more appear to Manoah and to his wife. Then Manoah knew that he was an angel of the LORD.
JUDG|13|22|And Manoah said unto his wife, We shall surely die, because we have seen God.
JUDG|13|23|But his wife said unto him, If the LORD were pleased to kill us, he would not have received a burnt offering and a meat offering at our hands, neither would he have showed us all these things, nor would as at this time have told us such things as these.
JUDG|13|24|And the woman bare a son, and called his name Samson: and the child grew, and the LORD blessed him.
JUDG|13|25|And the Spirit of the LORD began to move him at times in the camp of Dan between Zorah and Eshtaol.
JUDG|14|1|And Samson went down to Timnath, and saw a woman in Timnath of the daughters of the Philistines.
JUDG|14|2|And he came up, and told his father and his mother, and said, I have seen a woman in Timnath of the daughters of the Philistines: now therefore get her for me to wife.
JUDG|14|3|Then his father and his mother said unto him, Is there never a woman among the daughters of thy brethren, or among all my people, that thou goest to take a wife of the uncircumcised Philistines? And Samson said unto his father, Get her for me; for she pleaseth me well.
JUDG|14|4|But his father and his mother knew not that it was of the LORD, that he sought an occasion against the Philistines: for at that time the Philistines had dominion over Israel.
JUDG|14|5|Then went Samson down, and his father and his mother, to Timnath, and came to the vineyards of Timnath: and, behold, a young lion roared against him.
JUDG|14|6|And the Spirit of the LORD came mightily upon him, and he rent him as he would have rent a kid, and he had nothing in his hand: but he told not his father or his mother what he had done.
JUDG|14|7|And he went down, and talked with the woman; and she pleased Samson well.
JUDG|14|8|And after a time he returned to take her, and he turned aside to see the carcass of the lion: and, behold, there was a swarm of bees and honey in the carcass of the lion.
JUDG|14|9|And he took thereof in his hands, and went on eating, and came to his father and mother, and he gave them, and they did eat: but he told not them that he had taken the honey out of the carcass of the lion.
JUDG|14|10|So his father went down unto the woman: and Samson made there a feast; for so used the young men to do.
JUDG|14|11|And it came to pass, when they saw him, that they brought thirty companions to be with him.
JUDG|14|12|And Samson said unto them, I will now put forth a riddle unto you: if ye can certainly declare it me within the seven days of the feast, and find it out, then I will give you thirty sheets and thirty change of garments:
JUDG|14|13|But if ye cannot declare it me, then shall ye give me thirty sheets and thirty change of garments. And they said unto him, Put forth thy riddle, that we may hear it.
JUDG|14|14|And he said unto them, Out of the eater came forth meat, and out of the strong came forth sweetness. And they could not in three days expound the riddle.
JUDG|14|15|And it came to pass on the seventh day, that they said unto Samson's wife, Entice thy husband, that he may declare unto us the riddle, lest we burn thee and thy father's house with fire: have ye called us to take that we have? is it not so?
JUDG|14|16|And Samson's wife wept before him, and said, Thou dost but hate me, and lovest me not: thou hast put forth a riddle unto the children of my people, and hast not told it me. And he said unto her, Behold, I have not told it my father nor my mother, and shall I tell it thee?
JUDG|14|17|And she wept before him the seven days, while their feast lasted: and it came to pass on the seventh day, that he told her, because she lay sore upon him: and she told the riddle to the children of her people.
JUDG|14|18|And the men of the city said unto him on the seventh day before the sun went down, What is sweeter than honey? And what is stronger than a lion? and he said unto them, If ye had not plowed with my heifer, ye had not found out my riddle.
JUDG|14|19|And the Spirit of the LORD came upon him, and he went down to Ashkelon, and slew thirty men of them, and took their spoil, and gave change of garments unto them which expounded the riddle. And his anger was kindled, and he went up to his father's house.
JUDG|14|20|But Samson's wife was given to his companion, whom he had used as his friend.
JUDG|15|1|But it came to pass within a while after, in the time of wheat harvest, that Samson visited his wife with a kid; and he said, I will go in to my wife into the chamber. But her father would not suffer him to go in.
JUDG|15|2|And her father said, I verily thought that thou hadst utterly hated her; therefore I gave her to thy companion: is not her younger sister fairer than she? take her, I pray thee, instead of her.
JUDG|15|3|And Samson said concerning them, Now shall I be more blameless than the Philistines, though I do them a displeasure.
JUDG|15|4|And Samson went and caught three hundred foxes, and took firebrands, and turned tail to tail, and put a firebrand in the midst between two tails.
JUDG|15|5|And when he had set the brands on fire, he let them go into the standing corn of the Philistines, and burnt up both the shocks, and also the standing corn, with the vineyards and olives.
JUDG|15|6|Then the Philistines said, Who hath done this? And they answered, Samson, the son in law of the Timnite, because he had taken his wife, and given her to his companion. And the Philistines came up, and burnt her and her father with fire.
JUDG|15|7|And Samson said unto them, Though ye have done this, yet will I be avenged of you, and after that I will cease.
JUDG|15|8|And he smote them hip and thigh with a great slaughter: and he went down and dwelt in the top of the rock Etam.
JUDG|15|9|Then the Philistines went up, and pitched in Judah, and spread themselves in Lehi.
JUDG|15|10|And the men of Judah said, Why are ye come up against us? And they answered, To bind Samson are we come up, to do to him as he hath done to us.
JUDG|15|11|Then three thousand men of Judah went to the top of the rock Etam, and said to Samson, Knowest thou not that the Philistines are rulers over us? what is this that thou hast done unto us? And he said unto them, As they did unto me, so have I done unto them.
JUDG|15|12|And they said unto him, We are come down to bind thee, that we may deliver thee into the hand of the Philistines. And Samson said unto them, Swear unto me, that ye will not fall upon me yourselves.
JUDG|15|13|And they spake unto him, saying, No; but we will bind thee fast, and deliver thee into their hand: but surely we will not kill thee. And they bound him with two new cords, and brought him up from the rock.
JUDG|15|14|And when he came unto Lehi, the Philistines shouted against him: and the Spirit of the LORD came mightily upon him, and the cords that were upon his arms became as flax that was burnt with fire, and his bands loosed from off his hands.
JUDG|15|15|And he found a new jawbone of an ass, and put forth his hand, and took it, and slew a thousand men therewith.
JUDG|15|16|And Samson said, With the jawbone of an ass, heaps upon heaps, with the jaw of an ass have I slain a thousand men.
JUDG|15|17|And it came to pass, when he had made an end of speaking, that he cast away the jawbone out of his hand, and called that place Ramathlehi.
JUDG|15|18|And he was sore athirst, and called on the LORD, and said, Thou hast given this great deliverance into the hand of thy servant: and now shall I die for thirst, and fall into the hand of the uncircumcised?
JUDG|15|19|But God clave an hollow place that was in the jaw, and there came water thereout; and when he had drunk, his spirit came again, and he revived: wherefore he called the name thereof Enhakkore, which is in Lehi unto this day.
JUDG|15|20|And he judged Israel in the days of the Philistines twenty years.
JUDG|16|1|Then went Samson to Gaza, and saw there an harlot, and went in unto her.
JUDG|16|2|And it was told the Gazites, saying, Samson is come hither. And they compassed him in, and laid wait for him all night in the gate of the city, and were quiet all the night, saying, In the morning, when it is day, we shall kill him.
JUDG|16|3|And Samson lay till midnight, and arose at midnight, and took the doors of the gate of the city, and the two posts, and went away with them, bar and all, and put them upon his shoulders, and carried them up to the top of an hill that is before Hebron.
JUDG|16|4|And it came to pass afterward, that he loved a woman in the valley of Sorek, whose name was Delilah.
JUDG|16|5|And the lords of the Philistines came up unto her, and said unto her, Entice him, and see wherein his great strength lieth, and by what means we may prevail against him, that we may bind him to afflict him; and we will give thee every one of us eleven hundred pieces of silver.
JUDG|16|6|And Delilah said to Samson, Tell me, I pray thee, wherein thy great strength lieth, and wherewith thou mightest be bound to afflict thee.
JUDG|16|7|And Samson said unto her, If they bind me with seven green withes that were never dried, then shall I be weak, and be as another man.
JUDG|16|8|Then the lords of the Philistines brought up to her seven green withes which had not been dried, and she bound him with them.
JUDG|16|9|Now there were men lying in wait, abiding with her in the chamber. And she said unto him, The Philistines be upon thee, Samson. And he brake the withes, as a thread of tow is broken when it toucheth the fire. So his strength was not known.
JUDG|16|10|And Delilah said unto Samson, Behold, thou hast mocked me, and told me lies: now tell me, I pray thee, wherewith thou mightest be bound.
JUDG|16|11|And he said unto her, If they bind me fast with new ropes that never were occupied, then shall I be weak, and be as another man.
JUDG|16|12|Delilah therefore took new ropes, and bound him therewith, and said unto him, The Philistines be upon thee, Samson. And there were liers in wait abiding in the chamber. And he brake them from off his arms like a thread.
JUDG|16|13|And Delilah said unto Samson, Hitherto thou hast mocked me, and told me lies: tell me wherewith thou mightest be bound. And he said unto her, If thou weavest the seven locks of my head with the web.
JUDG|16|14|And she fastened it with the pin, and said unto him, The Philistines be upon thee, Samson. And he awaked out of his sleep, and went away with the pin of the beam, and with the web.
JUDG|16|15|And she said unto him, How canst thou say, I love thee, when thine heart is not with me? thou hast mocked me these three times, and hast not told me wherein thy great strength lieth.
JUDG|16|16|And it came to pass, when she pressed him daily with her words, and urged him, so that his soul was vexed unto death;
JUDG|16|17|That he told her all his heart, and said unto her, There hath not come a razor upon mine head; for I have been a Nazarite unto God from my mother's womb: if I be shaven, then my strength will go from me, and I shall become weak, and be like any other man.
JUDG|16|18|And when Delilah saw that he had told her all his heart, she sent and called for the lords of the Philistines, saying, Come up this once, for he hath showed me all his heart. Then the lords of the Philistines came up unto her, and brought money in their hand.
JUDG|16|19|And she made him sleep upon her knees; and she called for a man, and she caused him to shave off the seven locks of his head; and she began to afflict him, and his strength went from him.
JUDG|16|20|And she said, The Philistines be upon thee, Samson. And he awoke out of his sleep, and said, I will go out as at other times before, and shake myself. And he wist not that the LORD was departed from him.
JUDG|16|21|But the Philistines took him, and put out his eyes, and brought him down to Gaza, and bound him with fetters of brass; and he did grind in the prison house.
JUDG|16|22|Howbeit the hair of his head began to grow again after he was shaven.
JUDG|16|23|Then the lords of the Philistines gathered them together for to offer a great sacrifice unto Dagon their god, and to rejoice: for they said, Our god hath delivered Samson our enemy into our hand.
JUDG|16|24|And when the people saw him, they praised their god: for they said, Our god hath delivered into our hands our enemy, and the destroyer of our country, which slew many of us.
JUDG|16|25|And it came to pass, when their hearts were merry, that they said, Call for Samson, that he may make us sport. And they called for Samson out of the prison house; and he made them sport: and they set him between the pillars.
JUDG|16|26|And Samson said unto the lad that held him by the hand, Suffer me that I may feel the pillars whereupon the house standeth, that I may lean upon them.
JUDG|16|27|Now the house was full of men and women; and all the lords of the Philistines were there; and there were upon the roof about three thousand men and women, that beheld while Samson made sport.
JUDG|16|28|And Samson called unto the LORD, and said, O Lord God, remember me, I pray thee, and strengthen me, I pray thee, only this once, O God, that I may be at once avenged of the Philistines for my two eyes.
JUDG|16|29|And Samson took hold of the two middle pillars upon which the house stood, and on which it was borne up, of the one with his right hand, and of the other with his left.
JUDG|16|30|And Samson said, Let me die with the Philistines. And he bowed himself with all his might; and the house fell upon the lords, and upon all the people that were therein. So the dead which he slew at his death were more than they which he slew in his life.
JUDG|16|31|Then his brethren and all the house of his father came down, and took him, and brought him up, and buried him between Zorah and Eshtaol in the buryingplace of Manoah his father. And he judged Israel twenty years.
JUDG|17|1|And there was a man of mount Ephraim, whose name was Micah.
JUDG|17|2|And he said unto his mother, The eleven hundred shekels of silver that were taken from thee, about which thou cursedst, and spakest of also in mine ears, behold, the silver is with me; I took it. And his mother said, Blessed be thou of the LORD, my son.
JUDG|17|3|And when he had restored the eleven hundred shekels of silver to his mother, his mother said, I had wholly dedicated the silver unto the LORD from my hand for my son, to make a graven image and a molten image: now therefore I will restore it unto thee.
JUDG|17|4|Yet he restored the money unto his mother; and his mother took two hundred shekels of silver, and gave them to the founder, who made thereof a graven image and a molten image: and they were in the house of Micah.
JUDG|17|5|And the man Micah had an house of gods, and made an ephod, and teraphim, and consecrated one of his sons, who became his priest.
JUDG|17|6|In those days there was no king in Israel, but every man did that which was right in his own eyes.
JUDG|17|7|And there was a young man out of Bethlehemjudah of the family of Judah, who was a Levite, and he sojourned there.
JUDG|17|8|And the man departed out of the city from Bethlehemjudah to sojourn where he could find a place: and he came to mount Ephraim to the house of Micah, as he journeyed.
JUDG|17|9|And Micah said unto him, Whence comest thou? And he said unto him, I am a Levite of Bethlehemjudah, and I go to sojourn where I may find a place.
JUDG|17|10|And Micah said unto him, Dwell with me, and be unto me a father and a priest, and I will give thee ten shekels of silver by the year, and a suit of apparel, and thy victuals. So the Levite went in.
JUDG|17|11|And the Levite was content to dwell with the man; and the young man was unto him as one of his sons.
JUDG|17|12|And Micah consecrated the Levite; and the young man became his priest, and was in the house of Micah.
JUDG|17|13|Then said Micah, Now know I that the LORD will do me good, seeing I have a Levite to my priest.
JUDG|18|1|In those days there was no king in Israel: and in those days the tribe of the Danites sought them an inheritance to dwell in; for unto that day all their inheritance had not fallen unto them among the tribes of Israel.
JUDG|18|2|And the children of Dan sent of their family five men from their coasts, men of valor, from Zorah, and from Eshtaol, to spy out the land, and to search it; and they said unto them, Go, search the land: who when they came to mount Ephraim, to the house of Micah, they lodged there.
JUDG|18|3|When they were by the house of Micah, they knew the voice of the young man the Levite: and they turned in thither, and said unto him, Who brought thee hither? and what makest thou in this place? and what hast thou here?
JUDG|18|4|And he said unto them, Thus and thus dealeth Micah with me, and hath hired me, and I am his priest.
JUDG|18|5|And they said unto him, Ask counsel, we pray thee, of God, that we may know whether our way which we go shall be prosperous.
JUDG|18|6|And the priest said unto them, Go in peace: before the LORD is your way wherein ye go.
JUDG|18|7|Then the five men departed, and came to Laish, and saw the people that were therein, how they dwelt careless, after the manner of the Zidonians, quiet and secure; and there was no magistrate in the land, that might put them to shame in any thing; and they were far from the Zidonians, and had no business with any man.
JUDG|18|8|And they came unto their brethren to Zorah and Eshtaol: and their brethren said unto them, What say ye?
JUDG|18|9|And they said, Arise, that we may go up against them: for we have seen the land, and, behold, it is very good: and are ye still? be not slothful to go, and to enter to possess the land.
JUDG|18|10|When ye go, ye shall come unto a people secure, and to a large land: for God hath given it into your hands; a place where there is no want of any thing that is in the earth.
JUDG|18|11|And there went from thence of the family of the Danites, out of Zorah and out of Eshtaol, six hundred men appointed with weapons of war.
JUDG|18|12|And they went up, and pitched in Kirjathjearim, in Judah: wherefore they called that place Mahanehdan unto this day: behold, it is behind Kirjathjearim.
JUDG|18|13|And they passed thence unto mount Ephraim, and came unto the house of Micah.
JUDG|18|14|Then answered the five men that went to spy out the country of Laish, and said unto their brethren, Do ye know that there is in these houses an ephod, and teraphim, and a graven image, and a molten image? now therefore consider what ye have to do.
JUDG|18|15|And they turned thitherward, and came to the house of the young man the Levite, even unto the house of Micah, and saluted him.
JUDG|18|16|And the six hundred men appointed with their weapons of war, which were of the children of Dan, stood by the entering of the gate.
JUDG|18|17|And the five men that went to spy out the land went up, and came in thither, and took the graven image, and the ephod, and the teraphim, and the molten image: and the priest stood in the entering of the gate with the six hundred men that were appointed with weapons of war.
JUDG|18|18|And these went into Micah's house, and fetched the carved image, the ephod, and the teraphim, and the molten image. Then said the priest unto them, What do ye?
JUDG|18|19|And they said unto him, Hold thy peace, lay thine hand upon thy mouth, and go with us, and be to us a father and a priest: is it better for thee to be a priest unto the house of one man, or that thou be a priest unto a tribe and a family in Israel?
JUDG|18|20|And the priest's heart was glad, and he took the ephod, and the teraphim, and the graven image, and went in the midst of the people.
JUDG|18|21|So they turned and departed, and put the little ones and the cattle and the carriage before them.
JUDG|18|22|And when they were a good way from the house of Micah, the men that were in the houses near to Micah's house were gathered together, and overtook the children of Dan.
JUDG|18|23|And they cried unto the children of Dan. And they turned their faces, and said unto Micah, What aileth thee, that thou comest with such a company?
JUDG|18|24|And he said, Ye have taken away my gods which I made, and the priest, and ye are gone away: and what have I more? and what is this that ye say unto me, What aileth thee?
JUDG|18|25|And the children of Dan said unto him, Let not thy voice be heard among us, lest angry fellows run upon thee, and thou lose thy life, with the lives of thy household.
JUDG|18|26|And the children of Dan went their way: and when Micah saw that they were too strong for him, he turned and went back unto his house.
JUDG|18|27|And they took the things which Micah had made, and the priest which he had, and came unto Laish, unto a people that were at quiet and secure: and they smote them with the edge of the sword, and burnt the city with fire.
JUDG|18|28|And there was no deliverer, because it was far from Zidon, and they had no business with any man; and it was in the valley that lieth by Bethrehob. And they built a city, and dwelt therein.
JUDG|18|29|And they called the name of the city Dan, after the name of Dan their father, who was born unto Israel: howbeit the name of the city was Laish at the first.
JUDG|18|30|And the children of Dan set up the graven image: and Jonathan, the son of Gershom, the son of Manasseh, he and his sons were priests to the tribe of Dan until the day of the captivity of the land.
JUDG|18|31|And they set them up Micah's graven image, which he made, all the time that the house of God was in Shiloh.
JUDG|19|1|And it came to pass in those days, when there was no king in Israel, that there was a certain Levite sojourning on the side of mount Ephraim, who took to him a concubine out of Bethlehemjudah.
JUDG|19|2|And his concubine played the whore against him, and went away from him unto her father's house to Bethlehemjudah, and was there four whole months.
JUDG|19|3|And her husband arose, and went after her, to speak friendly unto her, and to bring her again, having his servant with him, and a couple of asses: and she brought him into her father's house: and when the father of the damsel saw him, he rejoiced to meet him.
JUDG|19|4|And his father in law, the damsel's father, retained him; and he abode with him three days: so they did eat and drink, and lodged there.
JUDG|19|5|And it came to pass on the fourth day, when they arose early in the morning, that he rose up to depart: and the damsel's father said unto his son in law, Comfort thine heart with a morsel of bread, and afterward go your way.
JUDG|19|6|And they sat down, and did eat and drink both of them together: for the damsel's father had said unto the man, Be content, I pray thee, and tarry all night, and let thine heart be merry.
JUDG|19|7|And when the man rose up to depart, his father in law urged him: therefore he lodged there again.
JUDG|19|8|And he arose early in the morning on the fifth day to depart; and the damsel's father said, Comfort thine heart, I pray thee. And they tarried until afternoon, and they did eat both of them.
JUDG|19|9|And when the man rose up to depart, he, and his concubine, and his servant, his father in law, the damsel's father, said unto him, Behold, now the day draweth toward evening, I pray you tarry all night: behold, the day groweth to an end, lodge here, that thine heart may be merry; and to morrow get you early on your way, that thou mayest go home.
JUDG|19|10|But the man would not tarry that night, but he rose up and departed, and came over against Jebus, which is Jerusalem; and there were with him two asses saddled, his concubine also was with him.
JUDG|19|11|And when they were by Jebus, the day was far spent; and the servant said unto his master, Come, I pray thee, and let us turn in into this city of the Jebusites, and lodge in it.
JUDG|19|12|And his master said unto him, We will not turn aside hither into the city of a stranger, that is not of the children of Israel; we will pass over to Gibeah.
JUDG|19|13|And he said unto his servant, Come, and let us draw near to one of these places to lodge all night, in Gibeah, or in Ramah.
JUDG|19|14|And they passed on and went their way; and the sun went down upon them when they were by Gibeah, which belongeth to Benjamin.
JUDG|19|15|And they turned aside thither, to go in and to lodge in Gibeah: and when he went in, he sat him down in a street of the city: for there was no man that took them into his house to lodging.
JUDG|19|16|And, behold, there came an old man from his work out of the field at even, which was also of mount Ephraim; and he sojourned in Gibeah: but the men of the place were Benjamites.
JUDG|19|17|And when he had lifted up his eyes, he saw a wayfaring man in the street of the city: and the old man said, Whither goest thou? and whence comest thou?
JUDG|19|18|And he said unto him, We are passing from Bethlehemjudah toward the side of mount Ephraim; from thence am I: and I went to Bethlehemjudah, but I am now going to the house of the LORD; and there is no man that receiveth me to house.
JUDG|19|19|Yet there is both straw and provender for our asses; and there is bread and wine also for me, and for thy handmaid, and for the young man which is with thy servants: there is no want of any thing.
JUDG|19|20|And the old man said, Peace be with thee; howsoever let all thy wants lie upon me; only lodge not in the street.
JUDG|19|21|So he brought him into his house, and gave provender unto the asses: and they washed their feet, and did eat and drink.
JUDG|19|22|Now as they were making their hearts merry, behold, the men of the city, certain sons of Belial, beset the house round about, and beat at the door, and spake to the master of the house, the old man, saying, Bring forth the man that came into thine house, that we may know him.
JUDG|19|23|And the man, the master of the house, went out unto them, and said unto them, Nay, my brethren, nay, I pray you, do not so wickedly; seeing that this man is come into mine house, do not this folly.
JUDG|19|24|Behold, here is my daughter a maiden, and his concubine; them I will bring out now, and humble ye them, and do with them what seemeth good unto you: but unto this man do not so vile a thing.
JUDG|19|25|But the men would not hearken to him: so the man took his concubine, and brought her forth unto them; and they knew her, and abused her all the night until the morning: and when the day began to spring, they let her go.
JUDG|19|26|Then came the woman in the dawning of the day, and fell down at the door of the man's house where her lord was, till it was light.
JUDG|19|27|And her lord rose up in the morning, and opened the doors of the house, and went out to go his way: and, behold, the woman his concubine was fallen down at the door of the house, and her hands were upon the threshold.
JUDG|19|28|And he said unto her, Up, and let us be going. But none answered. Then the man took her up upon an ass, and the man rose up, and gat him unto his place.
JUDG|19|29|And when he was come into his house, he took a knife, and laid hold on his concubine, and divided her, together with her bones, into twelve pieces, and sent her into all the coasts of Israel.
JUDG|19|30|And it was so, that all that saw it said, There was no such deed done nor seen from the day that the children of Israel came up out of the land of Egypt unto this day: consider of it, take advice, and speak your minds.
JUDG|20|1|Then all the children of Israel went out, and the congregation was gathered together as one man, from Dan even to Beersheba, with the land of Gilead, unto the LORD in Mizpeh.
JUDG|20|2|And the chief of all the people, even of all the tribes of Israel, presented themselves in the assembly of the people of God, four hundred thousand footmen that drew sword.
JUDG|20|3|(Now the children of Benjamin heard that the children of Israel were gone up to Mizpeh.) Then said the children of Israel, Tell us, how was this wickedness?
JUDG|20|4|And the Levite, the husband of the woman that was slain, answered and said, I came into Gibeah that belongeth to Benjamin, I and my concubine, to lodge.
JUDG|20|5|And the men of Gibeah rose against me, and beset the house round about upon me by night, and thought to have slain me: and my concubine have they forced, that she is dead.
JUDG|20|6|And I took my concubine, and cut her in pieces, and sent her throughout all the country of the inheritance of Israel: for they have committed lewdness and folly in Israel.
JUDG|20|7|Behold, ye are all children of Israel; give here your advice and counsel.
JUDG|20|8|And all the people arose as one man, saying, We will not any of us go to his tent, neither will we any of us turn into his house.
JUDG|20|9|But now this shall be the thing which we will do to Gibeah; we will go up by lot against it;
JUDG|20|10|And we will take ten men of an hundred throughout all the tribes of Israel, and an hundred of a thousand, and a thousand out of ten thousand, to fetch victual for the people, that they may do, when they come to Gibeah of Benjamin, according to all the folly that they have wrought in Israel.
JUDG|20|11|So all the men of Israel were gathered against the city, knit together as one man.
JUDG|20|12|And the tribes of Israel sent men through all the tribe of Benjamin, saying, What wickedness is this that is done among you?
JUDG|20|13|Now therefore deliver us the men, the children of Belial, which are in Gibeah, that we may put them to death, and put away evil from Israel. But the children of Benjamin would not hearken to the voice of their brethren the children of Israel.
JUDG|20|14|But the children of Benjamin gathered themselves together out of the cities unto Gibeah, to go out to battle against the children of Israel.
JUDG|20|15|And the children of Benjamin were numbered at that time out of the cities twenty and six thousand men that drew sword, beside the inhabitants of Gibeah, which were numbered seven hundred chosen men.
JUDG|20|16|Among all this people there were seven hundred chosen men lefthanded; every one could sling stones at an hair breadth, and not miss.
JUDG|20|17|And the men of Israel, beside Benjamin, were numbered four hundred thousand men that drew sword: all these were men of war.
JUDG|20|18|And the children of Israel arose, and went up to the house of God, and asked counsel of God, and said, Which of us shall go up first to the battle against the children of Benjamin? And the LORD said, Judah shall go up first.
JUDG|20|19|And the children of Israel rose up in the morning, and encamped against Gibeah.
JUDG|20|20|And the men of Israel went out to battle against Benjamin; and the men of Israel put themselves in array to fight against them at Gibeah.
JUDG|20|21|And the children of Benjamin came forth out of Gibeah, and destroyed down to the ground of the Israelites that day twenty and two thousand men.
JUDG|20|22|And the people the men of Israel encouraged themselves, and set their battle again in array in the place where they put themselves in array the first day.
JUDG|20|23|(And the children of Israel went up and wept before the LORD until even, and asked counsel of the LORD, saying, Shall I go up again to battle against the children of Benjamin my brother? And the LORD said, Go up against him.)
JUDG|20|24|And the children of Israel came near against the children of Benjamin the second day.
JUDG|20|25|And Benjamin went forth against them out of Gibeah the second day, and destroyed down to the ground of the children of Israel again eighteen thousand men; all these drew the sword.
JUDG|20|26|Then all the children of Israel, and all the people, went up, and came unto the house of God, and wept, and sat there before the LORD, and fasted that day until even, and offered burnt offerings and peace offerings before the LORD.
JUDG|20|27|And the children of Israel inquired of the LORD, (for the ark of the covenant of God was there in those days,
JUDG|20|28|And Phinehas, the son of Eleazar, the son of Aaron, stood before it in those days,) saying, Shall I yet again go out to battle against the children of Benjamin my brother, or shall I cease? And the LORD said, Go up; for to morrow I will deliver them into thine hand.
JUDG|20|29|And Israel set liers in wait round about Gibeah.
JUDG|20|30|And the children of Israel went up against the children of Benjamin on the third day, and put themselves in array against Gibeah, as at other times.
JUDG|20|31|And the children of Benjamin went out against the people, and were drawn away from the city; and they began to smite of the people, and kill, as at other times, in the highways, of which one goeth up to the house of God, and the other to Gibeah in the field, about thirty men of Israel.
JUDG|20|32|And the children of Benjamin said, They are smitten down before us, as at the first. But the children of Israel said, Let us flee, and draw them from the city unto the highways.
JUDG|20|33|And all the men of Israel rose up out of their place, and put themselves in array at Baaltamar: and the liers in wait of Israel came forth out of their places, even out of the meadows of Gibeah.
JUDG|20|34|And there came against Gibeah ten thousand chosen men out of all Israel, and the battle was sore: but they knew not that evil was near them.
JUDG|20|35|And the LORD smote Benjamin before Israel: and the children of Israel destroyed of the Benjamites that day twenty and five thousand and an hundred men: all these drew the sword.
JUDG|20|36|So the children of Benjamin saw that they were smitten: for the men of Israel gave place to the Benjamites, because they trusted unto the liers in wait which they had set beside Gibeah.
JUDG|20|37|And the liers in wait hasted, and rushed upon Gibeah; and the liers in wait drew themselves along, and smote all the city with the edge of the sword.
JUDG|20|38|Now there was an appointed sign between the men of Israel and the liers in wait, that they should make a great flame with smoke rise up out of the city.
JUDG|20|39|And when the men of Israel retired in the battle, Benjamin began to smite and kill of the men of Israel about thirty persons: for they said, Surely they are smitten down before us, as in the first battle.
JUDG|20|40|But when the flame began to arise up out of the city with a pillar of smoke, the Benjamites looked behind them, and, behold, the flame of the city ascended up to heaven.
JUDG|20|41|And when the men of Israel turned again, the men of Benjamin were amazed: for they saw that evil was come upon them.
JUDG|20|42|Therefore they turned their backs before the men of Israel unto the way of the wilderness; but the battle overtook them; and them which came out of the cities they destroyed in the midst of them.
JUDG|20|43|Thus they inclosed the Benjamites round about, and chased them, and trode them down with ease over against Gibeah toward the sunrising.
JUDG|20|44|And there fell of Benjamin eighteen thousand men; all these were men of valor.
JUDG|20|45|And they turned and fled toward the wilderness unto the rock of Rimmon: and they gleaned of them in the highways five thousand men; and pursued hard after them unto Gidom, and slew two thousand men of them.
JUDG|20|46|So that all which fell that day of Benjamin were twenty and five thousand men that drew the sword; all these were men of valor.
JUDG|20|47|But six hundred men turned and fled to the wilderness unto the rock Rimmon, and abode in the rock Rimmon four months.
JUDG|20|48|And the men of Israel turned again upon the children of Benjamin, and smote them with the edge of the sword, as well the men of every city, as the beast, and all that came to hand: also they set on fire all the cities that they came to.
JUDG|21|1|Now the men of Israel had sworn in Mizpeh, saying, There shall not any of us give his daughter unto Benjamin to wife.
JUDG|21|2|And the people came to the house of God, and abode there till even before God, and lifted up their voices, and wept sore;
JUDG|21|3|And said, O LORD God of Israel, why is this come to pass in Israel, that there should be to day one tribe lacking in Israel?
JUDG|21|4|And it came to pass on the morrow, that the people rose early, and built there an altar, and offered burnt offerings and peace offerings.
JUDG|21|5|And the children of Israel said, Who is there among all the tribes of Israel that came not up with the congregation unto the LORD? For they had made a great oath concerning him that came not up to the LORD to Mizpeh, saying, He shall surely be put to death.
JUDG|21|6|And the children of Israel repented them for Benjamin their brother, and said, There is one tribe cut off from Israel this day.
JUDG|21|7|How shall we do for wives for them that remain, seeing we have sworn by the LORD that we will not give them of our daughters to wives?
JUDG|21|8|And they said, What one is there of the tribes of Israel that came not up to Mizpeh to the LORD? And, behold, there came none to the camp from Jabeshgilead to the assembly.
JUDG|21|9|For the people were numbered, and, behold, there were none of the inhabitants of Jabeshgilead there.
JUDG|21|10|And the congregation sent thither twelve thousand men of the valiantest, and commanded them, saying, Go and smite the inhabitants of Jabeshgilead with the edge of the sword, with the women and the children.
JUDG|21|11|And this is the thing that ye shall do, Ye shall utterly destroy every male, and every woman that hath lain by man.
JUDG|21|12|And they found among the inhabitants of Jabeshgilead four hundred young virgins, that had known no man by lying with any male: and they brought them unto the camp to Shiloh, which is in the land of Canaan.
JUDG|21|13|And the whole congregation sent some to speak to the children of Benjamin that were in the rock Rimmon, and to call peaceably unto them.
JUDG|21|14|And Benjamin came again at that time; and they gave them wives which they had saved alive of the women of Jabeshgilead: and yet so they sufficed them not.
JUDG|21|15|And the people repented them for Benjamin, because that the LORD had made a breach in the tribes of Israel.
JUDG|21|16|Then the elders of the congregation said, How shall we do for wives for them that remain, seeing the women are destroyed out of Benjamin?
JUDG|21|17|And they said, There must be an inheritance for them that be escaped of Benjamin, that a tribe be not destroyed out of Israel.
JUDG|21|18|Howbeit we may not give them wives of our daughters: for the children of Israel have sworn, saying, Cursed be he that giveth a wife to Benjamin.
JUDG|21|19|Then they said, Behold, there is a feast of the LORD in Shiloh yearly in a place which is on the north side of Bethel, on the east side of the highway that goeth up from Bethel to Shechem, and on the south of Lebonah.
JUDG|21|20|Therefore they commanded the children of Benjamin, saying, Go and lie in wait in the vineyards;
JUDG|21|21|And see, and, behold, if the daughters of Shiloh come out to dance in dances, then come ye out of the vineyards, and catch you every man his wife of the daughters of Shiloh, and go to the land of Benjamin.
JUDG|21|22|And it shall be, when their fathers or their brethren come unto us to complain, that we will say unto them, Be favorable unto them for our sakes: because we reserved not to each man his wife in the war: for ye did not give unto them at this time, that ye should be guilty.
JUDG|21|23|And the children of Benjamin did so, and took them wives, according to their number, of them that danced, whom they caught: and they went and returned unto their inheritance, and repaired the cities, and dwelt in them.
JUDG|21|24|And the children of Israel departed thence at that time, every man to his tribe and to his family, and they went out from thence every man to his inheritance.
JUDG|21|25|In those days there was no king in Israel: every man did that which was right in his own eyes.
