HOS|1|1|当 乌西雅 、 约坦 、 亚哈斯 、 希西家 作 犹大 王， 约阿施 的儿子 耶罗波安 作 以色列 王的时候，耶和华的话临到 备利 的儿子 何西阿 。
HOS|1|2|耶和华初次向 何西阿 说话。耶和华对他说：“你去娶一个淫荡的女子为妻，收那从淫乱所生的儿女；因为这地行大淫乱，离弃耶和华。”
HOS|1|3|于是， 何西阿 去娶了 滴拉音 的女儿 歌篾 。她就怀孕，为 何西阿 生了一个儿子。
HOS|1|4|耶和华对 何西阿 说：“给他起名叫 耶斯列 ；因为再过片时，我要惩罚 耶户 家在 耶斯列 流人血的罪，也必终结 以色列 家的王朝。
HOS|1|5|到那日，我必在 耶斯列 平原折断 以色列 的弓。”
HOS|1|6|歌篾 又怀孕，生了一个女儿，耶和华对 何西阿 说：“给她起名叫 罗．路哈玛 ；因为我必不再怜悯 以色列 家，绝不赦免他们。
HOS|1|7|我却要怜悯 犹大 家，使他们靠耶和华－他们的上帝得救；我必不让他们靠弓、刀、战争、马匹与骑兵得救。”
HOS|1|8|歌篾 在 罗．路哈玛 断奶以后，又怀孕生了一个儿子。
HOS|1|9|耶和华说：“给他起名叫 罗．阿米 ；因为你们不是我的子民，我也不是你们的上帝 。”
HOS|1|10|然而， 以色列 的人数必多如海沙，不可量，不可数。从前在什么地方对他们说“你们不是我的子民”，将来就在那里称他们为“永生上帝的儿子”。
HOS|1|11|犹大 人和 以色列 人要一同聚集，为自己设立一个“头”，从这地上来，因为 耶斯列 的日子必为大日。
HOS|2|1|你们要称你们的众弟兄 为 阿米 ，称你们的众姊妹 为 路哈玛 。
HOS|2|2|要跟你们的母亲理论，理论， ─因为她不是我的妻子， 我也不是她的丈夫─ 叫她除掉脸上的淫相 和胸间的淫态，
HOS|2|3|免得我剥光她，使她赤身， 如刚出生的时候一样， 使她如旷野，如干旱之地， 干渴而死。
HOS|2|4|我必不怜悯她的儿女， 因为他们是从淫乱生的儿女。
HOS|2|5|他们的母亲行了淫乱， 怀他们的做了可羞耻的事； 因为她说：“我要跟随我所爱的， 我的饼、水、羊毛、麻、油、酒， 都是他们给的。”
HOS|2|6|因此，看哪，我要用荆棘堵塞她 的道， 筑墙挡住她， 使她找不着路；
HOS|2|7|以致她追随所爱的人，却追不上， 寻找他们，却寻不着， 就说：“我要回到前夫那里去， 因我那时比现在还好。”
HOS|2|8|她不知道是我给她五谷、新酒和新的油， 又加添她的金银； 他们却用来供奉 巴力 。
HOS|2|9|因此，我要在收割的日子收回我的五谷， 在当令的季节收回我的新酒， 我要夺回她用以遮体的羊毛和麻。
HOS|2|10|如今我必在她所爱的人眼前显露她的羞耻 ， 无人能救她脱离我的手。
HOS|2|11|我必使她的宴乐、节期、初一、安息日， 她一切的盛会都止息。
HOS|2|12|我要毁坏她的葡萄树和无花果树， 就是她所说“我所爱的给我为赏赐”的； 我要使它们变为荒林， 为野地的走兽所吞吃。
HOS|2|13|我要惩罚她素日给诸 巴力 烧香的罪； 那时她佩戴耳环和珠宝， 跟随她所爱的，却忘记我。 这是耶和华说的。
HOS|2|14|因此，看哪，我要诱导她，领她到旷野， 我要说动她的心。
HOS|2|15|在那里，我必赐她葡萄园， 又赐她 亚割谷 作为指望的门。 她必在那里回应， 像在年轻时从 埃及 地上来的时候一样。
HOS|2|16|那日你必称呼我 伊施 ，不再称呼我 巴力 。这是耶和华说的。
HOS|2|17|因为我必从她口中除掉诸 巴力 的名号，不再有人提这名号。
HOS|2|18|当那日，我必为我的百姓，与野地的走兽、天空的飞鸟和地上爬行的动物立约；又要在国中折断弓和刀，止息战争，使他们安然躺卧。
HOS|2|19|我必聘你永远归我为妻，以公义、公平、慈爱、怜悯聘你归我；
HOS|2|20|又以信实聘你归我，你就必认识耶和华。
HOS|2|21|耶和华说：那日我必应允， 我必应允天，天必应允地，
HOS|2|22|地必应允五谷、新酒和新的油； 这些都必应允在 耶斯列 身上。
HOS|2|23|我为自己必将她种在这地。 我必怜悯 罗．路哈玛 ； 对 罗．阿米 说： “你是我的子民”； 他必说：“我的上帝。”
HOS|3|1|耶和华又对我说：“你去爱那情人所爱却犯奸淫的妇人，正如耶和华爱那偏向别神、喜爱葡萄饼 的 以色列 人。”
HOS|3|2|于是我用十五舍客勒银子和一贺梅珥半大麦买她归我。
HOS|3|3|我对她说：“你当多日与我同住，不可行淫，不可归与别人，我对你也一样。”
HOS|3|4|因为 以色列 人必多日过着无君王，无领袖，无祭祀，无柱像，无以弗得，无家中神像的生活。
HOS|3|5|后来 以色列 人必归回 ，寻求耶和华─他们的上帝和他们的王 大卫 。在末后的日子，他们必敬畏耶和华，领受他的恩惠。
HOS|4|1|以色列 人哪，当听耶和华的话。 耶和华指控这地的居民， 因为在这地上无诚信， 无慈爱，无人认识上帝；
HOS|4|2|惟起誓、欺骗、杀害、 偷盗、奸淫、残暴、 流血又流血。
HOS|4|3|因此，这地悲哀， 其上的居民、野地的走兽、 天空的飞鸟都日趋衰微， 海中的鱼也必消灭。
HOS|4|4|然而，人都不必争辩，也不必指责。 你的百姓与抗拒祭司的人一样。
HOS|4|5|日间你必跌倒， 夜间先知也要与你一同跌倒； 我要灭绝你的母亲。
HOS|4|6|我的百姓因无知识而灭亡。 你抛弃知识， 我也必抛弃你， 使你不再作我的祭司。 你既忘了你上帝的律法， 我也必忘记你的儿女。
HOS|4|7|祭司越发增多，就越发得罪我； 我必使他们的荣耀变为羞辱。
HOS|4|8|他们吞吃我百姓的赎罪祭 ， 满心愿意我的子民犯罪。
HOS|4|9|将来百姓所受的， 祭司也必承受； 我必因他们所行的惩罚他们， 照他们所做的报应他们。
HOS|4|10|他们吃，却不得饱足； 行淫，却不繁衍； 因为他们离弃耶和华， 常行
HOS|4|11|淫乱。 酒和新酒夺去人的心。
HOS|4|12|我的百姓求问木头， 以为木杖能指示他们； 淫乱的心使他们失迷， 以致行淫离弃他们的上帝，
HOS|4|13|在各山顶献祭，在各高冈上烧香， 在橡树、杨树、大树之下， 因为那里树影美好。 所以，你们的女儿行淫， 你们的媳妇 犯奸淫。
HOS|4|14|我不因你们的女儿行淫 或你们的媳妇犯奸淫惩罚她们； 因为人自己转去与娼妓同居， 与神庙娼妓一同献祭。 这无知的百姓必致倾倒。
HOS|4|15|以色列 啊，你虽然行淫， 犹大 却不可犯罪； 不要往 吉甲 去， 不要上到 伯．亚文 ， 也不要指着永生的耶和华起誓。
HOS|4|16|以色列 倔强， 犹如倔强的母牛； 现在耶和华能牧放他们， 如在宽阔之地牧放羔羊吗？
HOS|4|17|以法莲 亲近偶像， 任凭他吧！
HOS|4|18|他们喝完了酒， 荒淫无度， 他们的官长甚爱羞耻的事。
HOS|4|19|风把他们卷在翅膀里， 他们必因所献的祭 蒙羞。
HOS|5|1|众祭司啊，要听这话！ 以色列 家啊，要留心听！ 王室啊，要侧耳而听！ 审判将临到你们， 因你们在 米斯巴 如罗网， 在 他泊山 如张开的网。
HOS|5|2|这些悖逆的人大行杀戮， 我要斥责他们众人。
HOS|5|3|至于我，我认识 以法莲 ， 以色列 不能向我隐藏。 以法莲 哪，现在你竟然行淫 ， 以色列 竟然被污辱。
HOS|5|4|他们所做的使他们不能归向上帝， 因有淫乱的心在他们里面； 他们不认识耶和华。
HOS|5|5|以色列 的骄傲使自己脸面无光 ； 以色列 和 以法莲 必因自己的罪孽跌倒， 犹大 也必与他们一同跌倒。
HOS|5|6|他们牵着牛羊去寻求耶和华， 却寻不着； 因他已转去离开他们。
HOS|5|7|他们不忠于耶和华， 生了私生子。 现在新月必吞灭他们和他们的地业。
HOS|5|8|你们当在 基比亚 吹角， 在 拉玛 吹号， 在 伯．亚文 发出警报； 便雅悯 哪，留意你的背后！
HOS|5|9|到了惩罚的日子， 以法莲 必变为废墟； 我在 以色列 众支派中，已指示将来必成的事。
HOS|5|10|犹大 的领袖如同挪移地界的人， 我必把我的愤怒如水倾倒在他们身上。
HOS|5|11|以法莲 因喜爱遵从荒谬的命令 就受欺压，在审判中被压碎。
HOS|5|12|我对 以法莲 竟如蛀虫， 向 犹大 家竟如朽烂。
HOS|5|13|以法莲 见自己有病， 犹大 见自己有伤， 以法莲 就前往 亚述 ， 差遣人去见大王 ； 他却不能医治你们， 不能治好你们的伤。
HOS|5|14|我必向 以法莲 如狮子， 向 犹大 家如少壮狮子。 我要撕裂，并且离去， 我必夺去，无人搭救。
HOS|5|15|我要去，我要回到原处， 等他们自觉有罪，寻求我的面； 急难时他们必切切寻求我。
HOS|6|1|来，我们归向耶和华吧！ 他撕裂我们，也必医治； 打伤我们，也必包扎。
HOS|6|2|过两天他必使我们苏醒， 第三天他必使我们兴起， 我们就在他面前得以存活。
HOS|6|3|我们要认识，要追求认识耶和华。 他如黎明必然出现， 他必临到我们像甘霖， 像滋润土地的春雨。
HOS|6|4|以法莲 哪，我可以向你怎样行呢？ 犹大 啊，我可以向你怎样做呢？ 因为你们的慈爱如同早晨的云雾， 又如速散的露水。
HOS|6|5|因此，我藉先知砍伐他们， 以我口中的话杀戮他们； 对你的审判 如光发出。
HOS|6|6|我喜爱慈爱 ，不喜爱祭物； 喜爱人认识上帝，胜于燔祭。
HOS|6|7|他们却如 亚当 背约， 在那里向我行诡诈。
HOS|6|8|基列 是作恶之人的城， 被血沾染。
HOS|6|9|成群的祭司如强盗埋伏等候， 在 示剑 的路上杀戮， 行了邪恶。
HOS|6|10|在 以色列 家我看见可憎的事， 在 以法莲 那里有淫行， 以色列 被污辱了。
HOS|6|11|犹大 啊，我使被掳之民归回的时候， 必有为你所预备的丰收。
HOS|7|1|我正要医治 以色列 的时候， 以法莲 的罪孽 和 撒玛利亚 的邪恶就显露出来。 他们行事虚谎， 内有贼人入侵， 外有群盗劫掠。
HOS|7|2|他们以为我不在意他们一切的恶行； 现在，他们所做的在我面前缠绕他们。
HOS|7|3|他们行恶使君王欢喜， 说谎使官长快乐。
HOS|7|4|他们全都犯奸淫， 如同烤热的火炉， 师傅在揉面到发面时 暂时停止煽火。
HOS|7|5|在我们君王宴乐的日子， 官长因酒的烈性而生病 ， 王与亵慢的人握手。
HOS|7|6|他们临近，心里如火炉一般， 他们等待，如烤饼的整夜睡觉， 到了早晨却如火焰熊熊。
HOS|7|7|他们全都热如火炉， 吞灭他们的审判官。 他们的君王都仆倒， 他们中间无一人求告我。
HOS|7|8|以法莲 混居在万民中 ， 以法莲 是没有翻过的饼。
HOS|7|9|外邦人消耗他的力量，他却不知道； 头发斑白，他也不觉得。
HOS|7|10|以色列 的骄傲使自己脸面无光。 他们虽遭遇这一切， 仍不归向耶和华－他们的上帝， 也不寻求他。
HOS|7|11|以法莲 好像鸽子愚蠢无知， 他们求告 埃及 ，投奔 亚述 。
HOS|7|12|他们去的时候，我要把我的网撒在他们身上； 我要捕获他们如同空中的鸟。 我必按他们会众所听到的 惩罚他们。
HOS|7|13|他们因离弃我，必定有祸； 因违背我，必遭毁灭。 我虽想要救赎他们，他们却向我说谎。
HOS|7|14|他们在床上呼号， 却不诚心哀求我； 他们为求五谷新酒而聚集 ， 却背叛我。
HOS|7|15|我虽管教他们，坚固他们的膀臂， 他们却图谋邪恶抗拒我。
HOS|7|16|他们归向，但不是归向至上者 ； 终究必如松弛的弓。 他们的领袖必因舌头的狂傲倒在刀下， 这在 埃及 地必成为人的笑柄。
HOS|8|1|你用口吹角吧！ 敌人如鹰攻打耶和华的家； 因为他们违背了我的约， 干犯了我的律法。
HOS|8|2|他们必呼求我： “我的上帝啊，我们 以色列 认识你了 。”
HOS|8|3|以色列 丢弃良善 ； 仇敌必追逼他。
HOS|8|4|他们立君王，并非出于我； 立官长，我却不知道。 他们用金银为自己制造偶像， 以致被剪除。
HOS|8|5|撒玛利亚 啊，耶和华已抛弃你的牛犊； 我的怒气向拜牛犊的人发作。 他们要到几时方能无罪呢？
HOS|8|6|因这牛犊是出于 以色列 ， 是匠人所造的， 并不是上帝。 撒玛利亚 的牛犊必被打碎。
HOS|8|7|他们所栽种的是风， 所收割的是暴风； 禾稼不长穗， 无以制成面粉； 即便制成， 外邦人也必吞吃它。
HOS|8|8|以色列 被吞吃， 如今在列国中像人所不喜爱的器皿。
HOS|8|9|他们投奔 亚述 如独行的野驴。 以法莲 雇用情人，
HOS|8|10|他们雇用列国； 如今我要聚集他们， 他们必因君王和官长所加的重担开始衰微 。
HOS|8|11|以法莲 为赎罪增添许多祭坛， 这些祭坛却使他犯罪。
HOS|8|12|我为他写了许多条 律法， 他却以为与他毫无关系。
HOS|8|13|他们献祭物作为给我的供物， 却自食其肉， 耶和华并不悦纳他们。 现在他必记起他们的罪孽， 惩罚他们的罪恶； 他们必返回 埃及 。
HOS|8|14|以色列 忘记造他的主，建造宫殿， 犹大 增添许多坚固的城； 我却要降火在他的城镇， 吞灭其堡垒。
HOS|9|1|以色列 啊，不要欢喜， 像 万民一样快乐； 因为你行淫离弃你的上帝， 喜爱各禾场上卖淫所得的赏金。
HOS|9|2|禾场和压酒池都不足以喂养他们， 它的新酒也必缺乏。
HOS|9|3|他们必不得住耶和华的地； 以法莲 却要返回 埃及 ， 在 亚述 吃不洁净的食物。
HOS|9|4|他们必不得向耶和华献浇酒祭， 所献的祭也不蒙悦纳。 他们的祭物如居丧者的食物， 凡吃的必使自己玷污； 因为他们的食物只为自己的口腹， 必不得入耶和华的殿。
HOS|9|5|到盛会的日子，在耶和华的节期， 你们要怎样行呢？
HOS|9|6|看哪，他们要逃避灾难； 埃及 人要收殓他们， 摩弗 人要埋葬他们。 蒺藜盘踞他们贵重的银器， 荆棘必占据他们的帐棚。
HOS|9|7|降罚的日子近了， 报应的时候已经来到。 以色列 必知道， 先知愚昧， 受灵感动的人狂妄， 皆因你多多作恶，大怀怨恨。
HOS|9|8|以法莲 替我的上帝守望； 至于先知，他所到之处都有捕鸟人的罗网， 在他上帝的家中也遭人怀恨。
HOS|9|9|他们深深败坏， 如在 基比亚 的日子一样。 耶和华必记起他们的罪孽， 惩罚他们的罪恶。
HOS|9|10|我发现 以色列 ， 如在旷野的葡萄； 我看见你们的祖先， 如春季无花果树上初熟的果子。 他们却来到 巴力．毗珥 ， 献上自己做羞耻的事， 成为可憎恶的， 与他们所爱的一样。
HOS|9|11|以法莲 ，他们的荣耀如鸟飞去， 必不生产，不怀胎，不成孕；
HOS|9|12|他们纵然将儿女养大， 我却要使他们丧子，一个也不留。 我离弃他们， 他们就有祸了。
HOS|9|13|我看 以法莲 如 推罗 栽于美地。 以法莲 却要将自己的儿女带出来， 交给行杀戮的人。
HOS|9|14|耶和华啊，求你加给他们， 加给他们什么呢？ 要使他们怀孕流产， 乳房枯干。
HOS|9|15|因他们在 吉甲 的一切恶事， 我在那里憎恶他们。 因他们所行的恶， 我必把他们赶出我的殿， 不再爱他们； 他们的领袖都是悖逆的。
HOS|9|16|以法莲 受击打， 其根枯干，不能结果， 即或生产， 我也要杀他们所生的爱子。
HOS|9|17|我的上帝必弃绝他们， 因为他们不听从他； 他们必飘流在列国中。
HOS|10|1|以色列 是茂盛的葡萄树， 结果繁多。 果子越多， 就越增添祭坛； 土地越肥美， 就越建造美丽的柱像。
HOS|10|2|他们心怀二意， 现今要定为有罪。 耶和华必拆毁他们的祭坛， 粉碎他们的柱像。
HOS|10|3|现在他们要说： “我们没有王； 因为我们不敬畏耶和华， 王又能为我们做什么呢？”
HOS|10|4|他们讲空话， 以假誓立约； 因此，惩罚如苦菜滋生 在田间的犁沟中。
HOS|10|5|撒玛利亚 的居民必因 伯．亚文 的牛犊惊恐； 它的百姓为它悲哀， 它的祭司为它战兢， 因为荣耀已经离开它。
HOS|10|6|人必将牛犊带到 亚述 ， 当作礼物献给大王。 以法莲 必蒙羞， 以色列 必因自己的计谋惭愧。
HOS|10|7|撒玛利亚 的王要灭亡， 如水面上的泡沫一般。
HOS|10|8|亚文 的丘坛， 以色列 犯罪的地方必毁坏， 荆棘和蒺藜必长在他们的祭坛上。 他们要向大山说：遮盖我们！ 向小山说：倒在我们身上！
HOS|10|9|以色列 啊， 你从 基比亚 的日子以来就时常犯罪， 他们仍停留在那里。 攻击罪孽之辈的战事岂不会临到 基比亚 吗？
HOS|10|10|我必随己意惩罚他们， 他们为双重的罪所缠； 万民必聚集攻击他们。
HOS|10|11|以法莲 是驯良的母牛犊，喜爱踹谷， 我要将轭套在它肥美的颈项上， 我要使 以法莲 被套住； 犹大 必耕田， 雅各 必耙地。
HOS|10|12|你们要为自己栽种公义， 收割慈爱。 你们要开垦荒地， 现今正是寻求耶和华的时候； 等他临到，公义必如雨降给你们。
HOS|10|13|你们耕种奸恶， 收割罪孽， 吃的是谎言的果实。 因你倚靠自己的行为， 仰赖你众多的勇士，
HOS|10|14|所以在你百姓中必掀起闹哄， 你一切的堡垒必被拆毁， 就如 沙勒幔 在争战的日子拆毁 伯．亚比勒 ， 将城中的母子一同摔死。
HOS|10|15|伯特利 啊，因你们的大恶， 你们必遭遇如此。 黎明来临， 以色列 的王必全然灭绝。
HOS|11|1|以色列 年幼的时候，我爱他， 就从 埃及 召我的儿子出来。
HOS|11|2|先知 越是呼唤他们， 他们越是远离 ， 向诸 巴力 献祭， 为雕刻的偶像烧香。
HOS|11|3|我曾教导 以法莲 行走， 我用膀臂 抱起他们， 他们却不知道是我医治他们。
HOS|11|4|我用慈绳爱索牵引他们； 我待他们如人松开牛两腮旁边的轭， 弯下身来喂养他们。
HOS|11|5|他们必不返回 埃及 地； 然而 亚述 人要作他们的王， 因他们不肯归向我。
HOS|11|6|刀剑必临到他们的城镇， 毁坏门闩，吞灭众人， 都因他们自己的计谋。
HOS|11|7|我的百姓偏要背离我， 他们虽向至高者呼求， 他却不抬举他们 。
HOS|11|8|以法莲 哪，我怎能舍弃你？ 以色列 啊，我怎能弃绝你？ 我怎能使你如 押玛 ？ 怎能使你如 洗扁 ？ 我回心转意， 我的怜悯燃了起来。
HOS|11|9|我必不发猛烈的怒气， 也不再毁灭 以法莲 。 因我是上帝，并非世人， 是你们中间的圣者； 我必不在怒中临到你们。
HOS|11|10|耶和华如狮子吼叫， 他的儿女必跟随他。 他一吼叫， 他们就从西方战兢而来。
HOS|11|11|他们必如雀鸟从 埃及 战兢而来， 又如鸽子从 亚述 地来到。 我必使他们住自己的房屋； 这是耶和华说的。
HOS|11|12|以法莲 用谎言围绕我， 以色列 家用诡计环绕我； 犹大 却仍与上帝同行 ， 向圣者忠心。
HOS|12|1|以法莲 以风为食物， 终日追逐东风， 增添虚谎和残暴， 与 亚述 立约， 也把油送到 埃及 。
HOS|12|2|耶和华指控 犹大 ， 要照 雅各 所行的惩罚他， 按他所做的报应他。
HOS|12|3|他在腹中抓住哥哥的脚跟， 壮年的时候与上帝角力，
HOS|12|4|他与天使角力，并且得胜。 他曾哀哭，恳求施恩。 在 伯特利 遇见耶和华， 耶和华在那里吩咐我们 ，
HOS|12|5|耶和华是万军之上帝， 耶和华是他可记念的名。
HOS|12|6|所以你当归向你的上帝， 谨守慈爱和公平， 常常等候你的上帝。
HOS|12|7|商人 手持诡诈的天平， 喜爱欺压。
HOS|12|8|以法莲 说： 我果然富有，得了财宝； 我所劳碌得来的一切 人必找不到我有什么可算为有罪的恶。
HOS|12|9|自从你出 埃及 地以来， 我就是耶和华－你的上帝； 我必使你再住帐棚， 如同节期的日子一样。
HOS|12|10|我已吩咐众先知， 又增加异象， 藉先知设比喻。
HOS|12|11|基列 没有罪孽吗？ 他们诚然是虚假的， 在 吉甲 献牛犊为祭； 他们的祭坛如同田间犁沟中的乱堆。
HOS|12|12|从前 雅各 逃到 亚兰 地， 以色列 为娶妻子工作， 为娶妻子而牧放。
HOS|12|13|后来耶和华藉先知领 以色列 从 埃及 上来， 也藉先知看顾他们。
HOS|12|14|然而 以法莲 大大惹动主怒， 他所流的血必归到他身上。 主必使他的羞辱归还给他。
HOS|13|1|从前 以法莲 说话，人都战兢， 他在 以色列 中居处高位； 但他因 巴力 犯罪就死了。
HOS|13|2|如今他们罪上加罪， 为自己铸造偶像， 凭自己的聪明用银子造偶像， 全都是匠人所制的。 论到它，有话说： 献祭的人都要亲吻牛犊。
HOS|13|3|因此，他们必如早晨的云雾， 又如速散的露水， 如被狂风吹离禾场的糠秕， 又如烟囱冒出的烟。
HOS|13|4|自从你出 埃及 地以来， 我就是耶和华－你的上帝； 除了我上帝以外，你不认识别的， 在我以外，并没有救主。
HOS|13|5|我曾在旷野， 就是那干旱之地认识你。
HOS|13|6|他们得到喂养，就饱足； 既得饱足，就心高气傲， 因而忘记了我。
HOS|13|7|因此我向他们如同狮子， 又如豹伏在道旁。
HOS|13|8|我如失去小熊的母熊，攻击他们， 撕裂他们的胸膛。 在那里我必如母狮吞吃他们， 如野兽撕开他们。
HOS|13|9|以色列 啊，你自取灭亡了 ， 因为我才是你的帮助。
HOS|13|10|现在，你的王在哪里呢？ 让他在你的各城中拯救你吧！ 你曾说“给我立君王和官长”， 那些治理你的又在哪里呢？
HOS|13|11|我在怒气中将王赐给你， 又在烈怒中将王废去。
HOS|13|12|以法莲 的罪孽被卷起来， 他的罪恶被收藏起来。
HOS|13|13|产妇的疼痛必临到他身上； 他是无智慧之子， 如同临盆时未出现的胎儿。
HOS|13|14|我必救赎他们脱离阴间， 救赎他们脱离死亡。 死亡啊，你的灾害在哪里？ 阴间哪，你的毁灭在哪里？ 怜悯必从我眼前消逝。
HOS|13|15|他在弟兄中虽然旺盛， 却有东风刮来， 就是耶和华的风从旷野上来。 他的泉源必干涸， 他的源头必枯竭， 这风必夺走他所积蓄的一切宝物。
HOS|13|16|撒玛利亚 要担当罪孽， 因为背叛自己的上帝。 他们必倒在刀下， 婴孩必被摔死， 孕妇必被剖开。
HOS|14|1|以色列 啊，你要归向耶和华－你的上帝， 你因自己的罪孽跌倒了。
HOS|14|2|当归向耶和华， 用言语向他说： “求你除尽罪孽，悦纳善行， 我们就用嘴唇的祭代替牛犊献上。
HOS|14|3|亚述 不能救我们， 我们不再骑马， 也不再对我们手所造的偶像说： ‘你是我们的上帝’； 孤儿在你那里得蒙怜悯。”
HOS|14|4|我必医治他们背道的病， 甘心爱他们， 因为我向他们所发的怒气已转消。
HOS|14|5|我必向 以色列 如甘露； 他必如百合花开放， 如 黎巴嫩 的树扎根。
HOS|14|6|他的嫩枝必延伸， 他的荣华如橄榄树， 香气如 黎巴嫩 的香柏树。
HOS|14|7|曾住在他荫下的必归回，使五谷生长 ， 他们要发旺如葡萄树， 他的名气 如 黎巴嫩 的酒。
HOS|14|8|以法莲 说： “我与偶像有何相干？” 我应允他，顾念他： 我如青翠的松树， 你的果实从我而来。
HOS|14|9|智慧人必明白这些事， 聪明人必知道这一切。 耶和华的道是正直的， 义人行在其中， 罪人却在其上跌倒。
