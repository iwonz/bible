HOS|1|1|The word of the LORD that came to Hosea son of Beeri during the reigns of Uzziah, Jotham, Ahaz and Hezekiah, kings of Judah, and during the reign of Jeroboam son of Jehoash king of Israel:
HOS|1|2|When the LORD began to speak through Hosea, the LORD said to him, "Go, take to yourself an adulterous wife and children of unfaithfulness, because the land is guilty of the vilest adultery in departing from the LORD."
HOS|1|3|So he married Gomer daughter of Diblaim, and she conceived and bore him a son.
HOS|1|4|Then the LORD said to Hosea, "Call him Jezreel, because I will soon punish the house of Jehu for the massacre at Jezreel, and I will put an end to the kingdom of Israel.
HOS|1|5|In that day I will break Israel's bow in the Valley of Jezreel."
HOS|1|6|Gomer conceived again and gave birth to a daughter. Then the LORD said to Hosea, "Call her Lo-Ruhamah, for I will no longer show love to the house of Israel, that I should at all forgive them.
HOS|1|7|Yet I will show love to the house of Judah; and I will save them-not by bow, sword or battle, or by horses and horsemen, but by the LORD their God."
HOS|1|8|After she had weaned Lo-Ruhamah, Gomer had another son.
HOS|1|9|Then the LORD said, "Call him Lo-Ammi, for you are not my people, and I am not your God.
HOS|1|10|"Yet the Israelites will be like the sand on the seashore, which cannot be measured or counted. In the place where it was said to them, 'You are not my people,' they will be called 'sons of the living God.'
HOS|1|11|The people of Judah and the people of Israel will be reunited, and they will appoint one leader and will come up out of the land, for great will be the day of Jezreel.
HOS|2|1|"Say of your brothers, 'My people,' and of your sisters, 'My loved one.'
HOS|2|2|"Rebuke your mother, rebuke her, for she is not my wife, and I am not her husband. Let her remove the adulterous look from her face and the unfaithfulness from between her breasts.
HOS|2|3|Otherwise I will strip her naked and make her as bare as on the day she was born; I will make her like a desert, turn her into a parched land, and slay her with thirst.
HOS|2|4|I will not show my love to her children, because they are the children of adultery.
HOS|2|5|Their mother has been unfaithful and has conceived them in disgrace. She said, 'I will go after my lovers, who give me my food and my water, my wool and my linen, my oil and my drink.'
HOS|2|6|Therefore I will block her path with thornbushes; I will wall her in so that she cannot find her way.
HOS|2|7|She will chase after her lovers but not catch them; she will look for them but not find them. Then she will say, 'I will go back to my husband as at first, for then I was better off than now.'
HOS|2|8|She has not acknowledged that I was the one who gave her the grain, the new wine and oil, who lavished on her the silver and gold- which they used for Baal.
HOS|2|9|"Therefore I will take away my grain when it ripens, and my new wine when it is ready. I will take back my wool and my linen, intended to cover her nakedness.
HOS|2|10|So now I will expose her lewdness before the eyes of her lovers; no one will take her out of my hands.
HOS|2|11|I will stop all her celebrations: her yearly festivals, her New Moons, her Sabbath days-all her appointed feasts.
HOS|2|12|I will ruin her vines and her fig trees, which she said were her pay from her lovers; I will make them a thicket, and wild animals will devour them.
HOS|2|13|I will punish her for the days she burned incense to the Baals; she decked herself with rings and jewelry, and went after her lovers, but me she forgot," declares the LORD.
HOS|2|14|"Therefore I am now going to allure her; I will lead her into the desert and speak tenderly to her.
HOS|2|15|There I will give her back her vineyards, and will make the Valley of Achor a door of hope. There she will sing as in the days of her youth, as in the day she came up out of Egypt.
HOS|2|16|"In that day," declares the LORD, "you will call me 'my husband'; you will no longer call me 'my master. '
HOS|2|17|I will remove the names of the Baals from her lips; no longer will their names be invoked.
HOS|2|18|In that day I will make a covenant for them with the beasts of the field and the birds of the air and the creatures that move along the ground. Bow and sword and battle I will abolish from the land, so that all may lie down in safety.
HOS|2|19|I will betroth you to me forever; I will betroth you in righteousness and justice, in love and compassion.
HOS|2|20|I will betroth you in faithfulness, and you will acknowledge the LORD.
HOS|2|21|"In that day I will respond," declares the LORD - "I will respond to the skies, and they will respond to the earth;
HOS|2|22|and the earth will respond to the grain, the new wine and oil, and they will respond to Jezreel.
HOS|2|23|I will plant her for myself in the land; I will show my love to the one I called 'Not my loved one. 'I will say to those called 'Not my people, You are my people'; and they will say, 'You are my God.'"
HOS|3|1|The LORD said to me, "Go, show your love to your wife again, though she is loved by another and is an adulteress. Love her as the LORD loves the Israelites, though they turn to other gods and love the sacred raisin cakes."
HOS|3|2|So I bought her for fifteen shekels of silver and about a homer and a lethek of barley.
HOS|3|3|Then I told her, "You are to live with me many days; you must not be a prostitute or be intimate with any man, and I will live with you."
HOS|3|4|For the Israelites will live many days without king or prince, without sacrifice or sacred stones, without ephod or idol.
HOS|3|5|Afterward the Israelites will return and seek the LORD their God and David their king. They will come trembling to the LORD and to his blessings in the last days.
HOS|4|1|Hear the word of the LORD, you Israelites, because the LORD has a charge to bring against you who live in the land: "There is no faithfulness, no love, no acknowledgment of God in the land.
HOS|4|2|There is only cursing, lying and murder, stealing and adultery; they break all bounds, and bloodshed follows bloodshed.
HOS|4|3|Because of this the land mourns, and all who live in it waste away; the beasts of the field and the birds of the air and the fish of the sea are dying.
HOS|4|4|"But let no man bring a charge, let no man accuse another, for your people are like those who bring charges against a priest.
HOS|4|5|You stumble day and night, and the prophets stumble with you. So I will destroy your mother-
HOS|4|6|my people are destroyed from lack of knowledge. "Because you have rejected knowledge, I also reject you as my priests; because you have ignored the law of your God, I also will ignore your children.
HOS|4|7|The more the priests increased, the more they sinned against me; they exchanged their Glory for something disgraceful.
HOS|4|8|They feed on the sins of my people and relish their wickedness.
HOS|4|9|And it will be: Like people, like priests. I will punish both of them for their ways and repay them for their deeds.
HOS|4|10|"They will eat but not have enough; they will engage in prostitution but not increase, because they have deserted the LORD to give themselves
HOS|4|11|to prostitution, to old wine and new, which take away the understanding
HOS|4|12|of my people. They consult a wooden idol and are answered by a stick of wood. A spirit of prostitution leads them astray; they are unfaithful to their God.
HOS|4|13|They sacrifice on the mountaintops and burn offerings on the hills, under oak, poplar and terebinth, where the shade is pleasant. Therefore your daughters turn to prostitution and your daughters-in-law to adultery.
HOS|4|14|"I will not punish your daughters when they turn to prostitution, nor your daughters-in-law when they commit adultery, because the men themselves consort with harlots and sacrifice with shrine prostitutes- a people without understanding will come to ruin!
HOS|4|15|"Though you commit adultery, O Israel, let not Judah become guilty. "Do not go to Gilgal; do not go up to Beth Aven. And do not swear, 'As surely as the LORD lives!'
HOS|4|16|The Israelites are stubborn, like a stubborn heifer. How then can the LORD pasture them like lambs in a meadow?
HOS|4|17|Ephraim is joined to idols; leave him alone!
HOS|4|18|Even when their drinks are gone, they continue their prostitution; their rulers dearly love shameful ways.
HOS|4|19|A whirlwind will sweep them away, and their sacrifices will bring them shame.
HOS|5|1|"Hear this, you priests! Pay attention, you Israelites! Listen, O royal house! This judgment is against you: You have been a snare at Mizpah, a net spread out on Tabor.
HOS|5|2|The rebels are deep in slaughter. I will discipline all of them.
HOS|5|3|I know all about Ephraim; Israel is not hidden from me. Ephraim, you have now turned to prostitution; Israel is corrupt.
HOS|5|4|"Their deeds do not permit them to return to their God. A spirit of prostitution is in their heart; they do not acknowledge the LORD.
HOS|5|5|Israel's arrogance testifies against them; the Israelites, even Ephraim, stumble in their sin; Judah also stumbles with them.
HOS|5|6|When they go with their flocks and herds to seek the LORD, they will not find him; he has withdrawn himself from them.
HOS|5|7|They are unfaithful to the LORD; they give birth to illegitimate children. Now their New Moon festivals will devour them and their fields.
HOS|5|8|"Sound the trumpet in Gibeah, the horn in Ramah. Raise the battle cry in Beth Aven; lead on, O Benjamin.
HOS|5|9|Ephraim will be laid waste on the day of reckoning. Among the tribes of Israel I proclaim what is certain.
HOS|5|10|Judah's leaders are like those who move boundary stones. I will pour out my wrath on them like a flood of water.
HOS|5|11|Ephraim is oppressed, trampled in judgment, intent on pursuing idols.
HOS|5|12|I am like a moth to Ephraim, like rot to the people of Judah.
HOS|5|13|"When Ephraim saw his sickness, and Judah his sores, then Ephraim turned to Assyria, and sent to the great king for help. But he is not able to cure you, not able to heal your sores.
HOS|5|14|For I will be like a lion to Ephraim, like a great lion to Judah. I will tear them to pieces and go away; I will carry them off, with no one to rescue them.
HOS|5|15|Then I will go back to my place until they admit their guilt. And they will seek my face; in their misery they will earnestly seek me."
HOS|6|1|"Come, let us return to the LORD. He has torn us to pieces but he will heal us; he has injured us but he will bind up our wounds.
HOS|6|2|After two days he will revive us; on the third day he will restore us, that we may live in his presence.
HOS|6|3|Let us acknowledge the LORD; let us press on to acknowledge him. As surely as the sun rises, he will appear; he will come to us like the winter rains, like the spring rains that water the earth."
HOS|6|4|"What can I do with you, Ephraim? What can I do with you, Judah? Your love is like the morning mist, like the early dew that disappears.
HOS|6|5|Therefore I cut you in pieces with my prophets, I killed you with the words of my mouth; my judgments flashed like lightning upon you.
HOS|6|6|For I desire mercy, not sacrifice, and acknowledgment of God rather than burnt offerings.
HOS|6|7|Like Adam, they have broken the covenant- they were unfaithful to me there.
HOS|6|8|Gilead is a city of wicked men, stained with footprints of blood.
HOS|6|9|As marauders lie in ambush for a man, so do bands of priests; they murder on the road to Shechem, committing shameful crimes.
HOS|6|10|I have seen a horrible thing in the house of Israel. There Ephraim is given to prostitution and Israel is defiled.
HOS|6|11|"Also for you, Judah, a harvest is appointed. "Whenever I would restore the fortunes of my people,
HOS|7|1|whenever I would heal Israel, the sins of Ephraim are exposed and the crimes of Samaria revealed. They practice deceit, thieves break into houses, bandits rob in the streets;
HOS|7|2|but they do not realize that I remember all their evil deeds. Their sins engulf them; they are always before me.
HOS|7|3|"They delight the king with their wickedness, the princes with their lies.
HOS|7|4|They are all adulterers, burning like an oven whose fire the baker need not stir from the kneading of the dough till it rises.
HOS|7|5|On the day of the festival of our king the princes become inflamed with wine, and he joins hands with the mockers.
HOS|7|6|Their hearts are like an oven; they approach him with intrigue. Their passion smolders all night; in the morning it blazes like a flaming fire.
HOS|7|7|All of them are hot as an oven; they devour their rulers. All their kings fall, and none of them calls on me.
HOS|7|8|"Ephraim mixes with the nations; Ephraim is a flat cake not turned over.
HOS|7|9|Foreigners sap his strength, but he does not realize it. His hair is sprinkled with gray, but he does not notice.
HOS|7|10|Israel's arrogance testifies against him, but despite all this he does not return to the LORD his God or search for him.
HOS|7|11|"Ephraim is like a dove, easily deceived and senseless- now calling to Egypt, now turning to Assyria.
HOS|7|12|When they go, I will throw my net over them; I will pull them down like birds of the air. When I hear them flocking together, I will catch them.
HOS|7|13|Woe to them, because they have strayed from me! Destruction to them, because they have rebelled against me! I long to redeem them but they speak lies against me.
HOS|7|14|They do not cry out to me from their hearts but wail upon their beds. They gather together for grain and new wine but turn away from me.
HOS|7|15|I trained them and strengthened them, but they plot evil against me.
HOS|7|16|They do not turn to the Most High; they are like a faulty bow. Their leaders will fall by the sword because of their insolent words. For this they will be ridiculed in the land of Egypt.
HOS|8|1|"Put the trumpet to your lips! An eagle is over the house of the LORD because the people have broken my covenant and rebelled against my law.
HOS|8|2|Israel cries out to me, 'O our God, we acknowledge you!'
HOS|8|3|But Israel has rejected what is good; an enemy will pursue him.
HOS|8|4|They set up kings without my consent; they choose princes without my approval. With their silver and gold they make idols for themselves to their own destruction.
HOS|8|5|Throw out your calf-idol, O Samaria! My anger burns against them. How long will they be incapable of purity?
HOS|8|6|They are from Israel! This calf-a craftsman has made it; it is not God. It will be broken in pieces, that calf of Samaria.
HOS|8|7|"They sow the wind and reap the whirlwind. The stalk has no head; it will produce no flour. Were it to yield grain, foreigners would swallow it up.
HOS|8|8|Israel is swallowed up; now she is among the nations like a worthless thing.
HOS|8|9|For they have gone up to Assyria like a wild donkey wandering alone. Ephraim has sold herself to lovers.
HOS|8|10|Although they have sold themselves among the nations, I will now gather them together. They will begin to waste away under the oppression of the mighty king.
HOS|8|11|"Though Ephraim built many altars for sin offerings, these have become altars for sinning.
HOS|8|12|I wrote for them the many things of my law, but they regarded them as something alien.
HOS|8|13|They offer sacrifices given to me and they eat the meat, but the LORD is not pleased with them. Now he will remember their wickedness and punish their sins: They will return to Egypt.
HOS|8|14|Israel has forgotten his Maker and built palaces; Judah has fortified many towns. But I will send fire upon their cities that will consume their fortresses."
HOS|9|1|Do not rejoice, O Israel; do not be jubilant like the other nations. For you have been unfaithful to your God; you love the wages of a prostitute at every threshing floor.
HOS|9|2|Threshing floors and winepresses will not feed the people; the new wine will fail them.
HOS|9|3|They will not remain in the LORD's land; Ephraim will return to Egypt and eat unclean food in Assyria.
HOS|9|4|They will not pour out wine offerings to the LORD, nor will their sacrifices please him. Such sacrifices will be to them like the bread of mourners; all who eat them will be unclean. This food will be for themselves; it will not come into the temple of the LORD.
HOS|9|5|What will you do on the day of your appointed feasts, on the festival days of the LORD?
HOS|9|6|Even if they escape from destruction, Egypt will gather them, and Memphis will bury them. Their treasures of silver will be taken over by briers, and thorns will overrun their tents.
HOS|9|7|The days of punishment are coming, the days of reckoning are at hand. Let Israel know this. Because your sins are so many and your hostility so great, the prophet is considered a fool, the inspired man a maniac.
HOS|9|8|The prophet, along with my God, is the watchman over Ephraim, yet snares await him on all his paths, and hostility in the house of his God.
HOS|9|9|They have sunk deep into corruption, as in the days of Gibeah. God will remember their wickedness and punish them for their sins.
HOS|9|10|"When I found Israel, it was like finding grapes in the desert; when I saw your fathers, it was like seeing the early fruit on the fig tree. But when they came to Baal Peor, they consecrated themselves to that shameful idol and became as vile as the thing they loved.
HOS|9|11|Ephraim's glory will fly away like a bird- no birth, no pregnancy, no conception.
HOS|9|12|Even if they rear children, I will bereave them of every one. Woe to them when I turn away from them!
HOS|9|13|I have seen Ephraim, like Tyre, planted in a pleasant place. But Ephraim will bring out their children to the slayer."
HOS|9|14|Give them, O LORD - what will you give them? Give them wombs that miscarry and breasts that are dry.
HOS|9|15|"Because of all their wickedness in Gilgal, I hated them there. Because of their sinful deeds, I will drive them out of my house. I will no longer love them; all their leaders are rebellious.
HOS|9|16|Ephraim is blighted, their root is withered, they yield no fruit. Even if they bear children, I will slay their cherished offspring."
HOS|9|17|My God will reject them because they have not obeyed him; they will be wanderers among the nations.
HOS|10|1|Israel was a spreading vine; he brought forth fruit for himself. As his fruit increased, he built more altars; as his land prospered, he adorned his sacred stones.
HOS|10|2|Their heart is deceitful, and now they must bear their guilt. The LORD will demolish their altars and destroy their sacred stones.
HOS|10|3|Then they will say, "We have no king because we did not revere the LORD. But even if we had a king, what could he do for us?"
HOS|10|4|They make many promises, take false oaths and make agreements; therefore lawsuits spring up like poisonous weeds in a plowed field.
HOS|10|5|The people who live in Samaria fear for the calf-idol of Beth Aven. Its people will mourn over it, and so will its idolatrous priests, those who had rejoiced over its splendor, because it is taken from them into exile.
HOS|10|6|It will be carried to Assyria as tribute for the great king. Ephraim will be disgraced; Israel will be ashamed of its wooden idols.
HOS|10|7|Samaria and its king will float away like a twig on the surface of the waters.
HOS|10|8|The high places of wickedness will be destroyed- it is the sin of Israel. Thorns and thistles will grow up and cover their altars. Then they will say to the mountains, "Cover us!" and to the hills, "Fall on us!"
HOS|10|9|"Since the days of Gibeah, you have sinned, O Israel, and there you have remained. Did not war overtake the evildoers in Gibeah?
HOS|10|10|When I please, I will punish them; nations will be gathered against them to put them in bonds for their double sin.
HOS|10|11|Ephraim is a trained heifer that loves to thresh; so I will put a yoke on her fair neck. I will drive Ephraim, Judah must plow, and Jacob must break up the ground.
HOS|10|12|Sow for yourselves righteousness, reap the fruit of unfailing love, and break up your unplowed ground; for it is time to seek the LORD, until he comes and showers righteousness on you.
HOS|10|13|But you have planted wickedness, you have reaped evil, you have eaten the fruit of deception. Because you have depended on your own strength and on your many warriors,
HOS|10|14|the roar of battle will rise against your people, so that all your fortresses will be devastated- as Shalman devastated Beth Arbel on the day of battle, when mothers were dashed to the ground with their children.
HOS|10|15|Thus will it happen to you, O Bethel, because your wickedness is great. When that day dawns, the king of Israel will be completely destroyed.
HOS|11|1|"When Israel was a child, I loved him, and out of Egypt I called my son.
HOS|11|2|But the more I called Israel, the further they went from me. They sacrificed to the Baals and they burned incense to images.
HOS|11|3|It was I who taught Ephraim to walk, taking them by the arms; but they did not realize it was I who healed them.
HOS|11|4|I led them with cords of human kindness, with ties of love; I lifted the yoke from their neck and bent down to feed them.
HOS|11|5|"Will they not return to Egypt and will not Assyria rule over them because they refuse to repent?
HOS|11|6|Swords will flash in their cities, will destroy the bars of their gates and put an end to their plans.
HOS|11|7|My people are determined to turn from me. Even if they call to the Most High, he will by no means exalt them.
HOS|11|8|"How can I give you up, Ephraim? How can I hand you over, Israel? How can I treat you like Admah? How can I make you like Zeboiim? My heart is changed within me; all my compassion is aroused.
HOS|11|9|I will not carry out my fierce anger, nor will I turn and devastate Ephraim. For I am God, and not man- the Holy One among you. I will not come in wrath.
HOS|11|10|They will follow the LORD; he will roar like a lion. When he roars, his children will come trembling from the west.
HOS|11|11|They will come trembling like birds from Egypt, like doves from Assyria. I will settle them in their homes," declares the LORD.
HOS|11|12|Ephraim has surrounded me with lies, the house of Israel with deceit. And Judah is unruly against God, even against the faithful Holy One.
HOS|12|1|Ephraim feeds on the wind; he pursues the east wind all day and multiplies lies and violence. He makes a treaty with Assyria and sends olive oil to Egypt.
HOS|12|2|The LORD has a charge to bring against Judah; he will punish Jacob according to his ways and repay him according to his deeds.
HOS|12|3|In the womb he grasped his brother's heel; as a man he struggled with God.
HOS|12|4|He struggled with the angel and overcame him; he wept and begged for his favor. He found him at Bethel and talked with him there-
HOS|12|5|the LORD God Almighty, the LORD is his name of renown!
HOS|12|6|But you must return to your God; maintain love and justice, and wait for your God always.
HOS|12|7|The merchant uses dishonest scales; he loves to defraud.
HOS|12|8|Ephraim boasts, "I am very rich; I have become wealthy. With all my wealth they will not find in me any iniquity or sin."
HOS|12|9|"I am the LORD your God, who brought you out of Egypt; I will make you live in tents again, as in the days of your appointed feasts.
HOS|12|10|I spoke to the prophets, gave them many visions and told parables through them."
HOS|12|11|Is Gilead wicked? Its people are worthless! Do they sacrifice bulls in Gilgal? Their altars will be like piles of stones on a plowed field.
HOS|12|12|Jacob fled to the country of Aram; Israel served to get a wife, and to pay for her he tended sheep.
HOS|12|13|The LORD used a prophet to bring Israel up from Egypt, by a prophet he cared for him.
HOS|12|14|But Ephraim has bitterly provoked him to anger; his Lord will leave upon him the guilt of his bloodshed and will repay him for his contempt.
HOS|13|1|When Ephraim spoke, men trembled; he was exalted in Israel. But he became guilty of Baal worship and died.
HOS|13|2|Now they sin more and more; they make idols for themselves from their silver, cleverly fashioned images, all of them the work of craftsmen. It is said of these people, "They offer human sacrifice and kiss the calf-idols."
HOS|13|3|Therefore they will be like the morning mist, like the early dew that disappears, like chaff swirling from a threshing floor, like smoke escaping through a window.
HOS|13|4|"But I am the LORD your God, who brought you out of Egypt. You shall acknowledge no God but me, no Savior except me.
HOS|13|5|I cared for you in the desert, in the land of burning heat.
HOS|13|6|When I fed them, they were satisfied; when they were satisfied, they became proud; then they forgot me.
HOS|13|7|So I will come upon them like a lion, like a leopard I will lurk by the path.
HOS|13|8|Like a bear robbed of her cubs, I will attack them and rip them open. Like a lion I will devour them; a wild animal will tear them apart.
HOS|13|9|"You are destroyed, O Israel, because you are against me, against your helper.
HOS|13|10|Where is your king, that he may save you? Where are your rulers in all your towns, of whom you said, 'Give me a king and princes'?
HOS|13|11|So in my anger I gave you a king, and in my wrath I took him away.
HOS|13|12|The guilt of Ephraim is stored up, his sins are kept on record.
HOS|13|13|Pains as of a woman in childbirth come to him, but he is a child without wisdom; when the time arrives, he does not come to the opening of the womb.
HOS|13|14|"I will ransom them from the power of the grave; I will redeem them from death. Where, O death, are your plagues? Where, O grave, is your destruction? "I will have no compassion,
HOS|13|15|even though he thrives among his brothers. An east wind from the LORD will come, blowing in from the desert; his spring will fail and his well dry up. His storehouse will be plundered of all its treasures.
HOS|13|16|The people of Samaria must bear their guilt, because they have rebelled against their God. They will fall by the sword; their little ones will be dashed to the ground, their pregnant women ripped open."
HOS|14|1|Return, O Israel, to the LORD your God. Your sins have been your downfall!
HOS|14|2|Take words with you and return to the LORD. Say to him: "Forgive all our sins and receive us graciously, that we may offer the fruit of our lips.
HOS|14|3|Assyria cannot save us; we will not mount war-horses. We will never again say 'Our gods' to what our own hands have made, for in you the fatherless find compassion."
HOS|14|4|"I will heal their waywardness and love them freely, for my anger has turned away from them.
HOS|14|5|I will be like the dew to Israel; he will blossom like a lily. Like a cedar of Lebanon he will send down his roots;
HOS|14|6|his young shoots will grow. His splendor will be like an olive tree, his fragrance like a cedar of Lebanon.
HOS|14|7|Men will dwell again in his shade. He will flourish like the grain. He will blossom like a vine, and his fame will be like the wine from Lebanon.
HOS|14|8|O Ephraim, what more have I to do with idols? I will answer him and care for him. I am like a green pine tree; your fruitfulness comes from me."
HOS|14|9|Who is wise? He will realize these things. Who is discerning? He will understand them. The ways of the LORD are right; the righteous walk in them, but the rebellious stumble in them.
