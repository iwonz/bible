JER|1|1|这些是 便雅悯 地 亚拿突城 的祭司， 希勒家 的儿子 耶利米 的话。
JER|1|2|亚们 的儿子 犹大 王 约西亚 在位第十三年，耶和华的话临到 耶利米 。
JER|1|3|从 约西亚 的儿子 犹大 王 约雅敬 在位的时候，直到 约西亚 的儿子 犹大 王 西底家 在位的末年，就是第十一年五月间 耶路撒冷 被掳时，耶和华的话也常临到 耶利米 。
JER|1|4|耶利米 说，耶和华的话临到我，说：
JER|1|5|“我尚未将你造在母腹中，就已认识你； 你未出母胎，我已将你分别为圣， 派你作列国的先知。”
JER|1|6|我就说：“唉，主耶和华！看哪，我不知道怎么说，因为我年轻。”
JER|1|7|耶和华对我说： “不要说：‘我年轻’， 因为我差遣你到谁那里去，你都要去； 我吩咐你说什么话，你都要说。
JER|1|8|你不要怕他们， 因为我与你同在，要拯救你。 这是耶和华说的。”
JER|1|9|于是耶和华伸手按住我的口， 对我说： “看哪，我已将我的话放在你口中。
JER|1|10|我今日立你在列邦列国之上， 为要拔出，拆毁，毁坏，倾覆， 又要建立，栽植。”
JER|1|11|耶和华的话临到我，说：“ 耶利米 ，你看见什么？”我说：“我看见一根杏树枝。”
JER|1|12|耶和华对我说：“你看得不错；因为我要看守 我的话，使它实现。”
JER|1|13|耶和华的话第二次临到我，说：“你看见什么？”我说：“我看见一个水烧开的锅，从北而倾。”
JER|1|14|耶和华对我说：“必有灾祸从北方发出，临到这地所有的居民。
JER|1|15|看哪，我要召北方列国的万族。这是耶和华说的。他们要来，各安宝座在 耶路撒冷 的城门口，周围攻击城墙，又要攻击 犹大 的一切城镇。
JER|1|16|这百姓离弃我，向别神烧香，跪拜自己手所造的，我要针对这一切恶行，向他们宣读我的判决。
JER|1|17|所以你当束腰，起来，将我所吩咐你的一切话都告诉他们；不要因他们惊惶，免得我使你在他们面前惊惶。
JER|1|18|看哪，我今日使你成为坚城、铁柱、铜墙，对抗全地和 犹大 的君王、官长、祭司，并这地的百姓。
JER|1|19|他们要攻击你，却不能胜过你，因为我与你同在，要拯救你。这是耶和华说的。”
JER|2|1|耶和华的话临到我，说：
JER|2|2|“你去向 耶路撒冷 居民的耳朵呼喊说，耶和华如此说： ‘你年轻时的恩爱， 新婚时的爱情， 你怎样在旷野， 在未耕种之地跟随我， 我都记得。
JER|2|3|那时 以色列 归耶和华为圣， 作为他初熟的土产； 凡吞吃它的必算为有罪， 灾祸必临到他们。 这是耶和华说的。’”
JER|2|4|雅各 家， 以色列 家的各族啊，当听耶和华的话，
JER|2|5|耶和华如此说： “你们的祖先看我有什么错处， 竟远离我，随从那虚无的神明 ， 自己成为虚无呢？
JER|2|6|他们并不问： ‘那领我们从 埃及 地上来， 引导我们走过旷野、沙漠有坑洞之地， 走过干旱死荫、无人经过、 无人居住之地的耶和华在哪里呢？’
JER|2|7|我领你们进入肥沃之地， 使你们得吃其中的果子和美物； 你们进入时，却使我的地玷污， 使我的产业成为可憎恶的。
JER|2|8|祭司从来不问：‘耶和华在哪里呢？’ 传讲律法的不认识我， 官长违背我， 先知藉 巴力 说预言， 随从无益的东西。”
JER|2|9|“我因此必与你们争辩， 也与你们的子孙争辩。 这是耶和华说的。
JER|2|10|你们且渡到 基提 海岛察看， 派人往 基达 去留心查考， 看可曾有过这样的事。
JER|2|11|岂有一国换了它的神明吗？ 其实那不是神明！ 但我的百姓将他们的荣耀换了那无益的东西。
JER|2|12|诸天哪，要因此震惊， 颤栗，极其凄凉！ 这是耶和华说的。
JER|2|13|因为我的百姓做了两件恶事： 离弃我这活水的泉源； 又为自己凿出水池， 却是破裂不能储水的池子。”
JER|2|14|“ 以色列 是仆人吗？ 是家中生的奴仆吗？ 为何成为掠物呢？
JER|2|15|少壮狮子向它咆哮，大声吼叫， 使它的地荒芜； 城镇烧毁，无人居住。
JER|2|16|挪弗 人和 答比匿 人打破你的头颅。
JER|2|17|这不是你自己招惹的吗？ 不是因耶和华－你上帝引导你行路时， 你离弃了他吗？
JER|2|18|现今你为何在 埃及 路上喝 西曷河 的水呢？ 为何在 亚述 路上喝 大河 的水呢？
JER|2|19|你自己的恶必惩治你， 你背道的事必责罚你。 由此可知可见，你离弃耶和华－你的上帝， 不存敬畏我的心， 实为恶事，为苦事； 这是万军之主耶和华说的。”
JER|2|20|“你 在古时折断你的轭，解开你的绳索， 说：‘我必不事奉耶和华 。’ 你在各高冈上、各青翠的树下屈身行淫。
JER|2|21|然而，我栽种你为上等的葡萄树， 全用纯正的种子； 你怎么向我变为外邦葡萄树的坏枝子呢？
JER|2|22|你虽用碱、多用皂荚清洗， 你罪孽的痕迹仍显在我面前。 这是主耶和华说的。
JER|2|23|你怎能说： ‘我没有玷污，没有随从 巴力 ’？ 看看你在谷中所做的，思想你自己的所作所为； 你是快行的独峰驼，狂奔乱闯。
JER|2|24|你是野驴，习惯旷野， 欲心发动时就呼吸急促， 发情时谁能使它转回呢？ 凡寻找它的必不费力， 在它的季节必能寻见它。
JER|2|25|你不要弄到赤足而行， 喉咙干渴。 你却说：‘没有用的， 我喜爱陌生人， 我必随从他们。’”
JER|2|26|“贼被捉拿，怎样羞愧， 以色列 家和他们的君王、官长、 祭司、先知也都照样羞愧。
JER|2|27|他们向木头说：‘你是我的父’； 向石头说：‘你是生我的。’ 他们以背向我， 不肯以面向我； 及至遭遇患难时却说： ‘起来拯救我们吧！’
JER|2|28|你为自己做的神明在哪里呢？ 你遭遇患难的时候， 让它们起来拯救你吧！ 犹大 啊，你神明的数目与你城的数目相等。
JER|2|29|“你们为何与我争辩呢？ 你们都违背了我。 这是耶和华说的。
JER|2|30|我责打你们的儿女是徒然的， 他们不受管教。 你们自己的刀吞灭你们的先知， 好像残害人的狮子。
JER|2|31|这世代的人哪， 你们要留意耶和华的话。 我向 以色列 岂是旷野， 或幽暗之地呢？ 我的百姓为何说： ‘我们脱离约束，不再归向你了’？
JER|2|32|少女岂能忘记她的妆饰呢？ 新娘岂能忘记她的美衣呢？ 我的百姓却在无数的日子里忘记了我！
JER|2|33|“你竟然如此精于求爱之道， 可把你的门径教邪恶的女人！
JER|2|34|你衣服的边上有无辜贫穷人的血， 其实你并未发现他们挖洞进屋偷窃 。 虽有这一切的事 ，
JER|2|35|你还说：‘我无辜； 耶和华的怒气必定转离我了。’ 看哪，我必审问你； 因你自己说：‘我没有犯罪。’
JER|2|36|你为何东奔西跑改变你的道路呢？ 你必因 埃及 蒙羞， 像从前因 亚述 蒙羞一样。
JER|2|37|你也必两手抱头离开这里； 因为耶和华已经弃绝你所倚靠的， 你不能因他们而得顺利。”
JER|3|1|耶和华说 ：“人若休妻， 妻离他而去，做了别人的妻子， 前夫岂能再回到她那里呢？ 那地岂不是大大污秽了吗？ 但你和许多情郎行淫， 还是可以回到我这里。 这是耶和华说的。
JER|3|2|你举目向光秃的高地观看， 何处没有你的淫行呢？ 你坐在道路旁等候， 好像 阿拉伯 人在旷野埋伏， 你的淫行和邪恶使全地污秽了。
JER|3|3|因此甘霖停止， 春雨不降。 你还是一副娼妓之脸， 不顾羞耻。
JER|3|4|你不是才向我呼叫说： ‘我父啊，你是我年轻时的密友，
JER|3|5|人岂永远怀恨，长久存怒吗？’ 看哪，你虽这样说，还是竭尽所能去行恶。”
JER|3|6|约西亚 王在位的时候，耶和华对我说：“你看见背道的 以色列 所做的吗？她上到各高山，在各青翠的树下行淫。
JER|3|7|我说：‘她行这些事以后会回转归向我’，她却不回转。她奸诈的妹妹 犹大 也看见了。
JER|3|8|我看见背道的 以色列 行淫，我为这缘故给她休书休了她，她奸诈的妹妹 犹大 还不惧怕，也去行淫。
JER|3|9|因 以色列 轻忽了她的淫乱，与石头和木头行奸淫 ，她和这地就都污秽了 。
JER|3|10|虽有这一切的事，她奸诈的妹妹 犹大 还不一心归向我，不过是假意归我。这是耶和华说的。”
JER|3|11|耶和华对我说：“背道的 以色列 比奸诈的 犹大 还显为义。
JER|3|12|你去向北方宣告这些话，说： ‘背道的 以色列 啊，回来吧！ 这是耶和华说的。 我必不怒目看你们， 因为我是慈爱的， 这是耶和华说的。 我必不永远怀怒；
JER|3|13|只要你承认你的罪孽， 就是违背耶和华－你的上帝， 在各青翠的树下追逐外族的神明 ， 没有听从我的话。 这是耶和华说的。
JER|3|14|背道的儿女啊，回来吧！ 这是耶和华说的。 因为我作你们的丈夫， 要将你们从一城取一人， 从一族取两人，带到 锡安 。
JER|3|15|“‘我必将合我心意的牧者赏赐给你们，他们要以知识和智慧牧养你们。
JER|3|16|你们在国中生养众多的时候，那些日子，人必不再提说耶和华的约柜，不追想，不记念，不觉缺少，也不再制造。这是耶和华说的。
JER|3|17|那时，人必称 耶路撒冷 为耶和华的宝座；万国聚集在那里，为耶和华的名来到 耶路撒冷 ，他们必不再随从自己顽梗的恶心行事。
JER|3|18|当那些日子， 犹大 家要和 以色列 家同行，从北方之地一同来到我所赐给你们祖先为业之地。’”
JER|3|19|我说，我多么乐意把你列在儿女之中， 赐给你美地， 就是万国中最美的产业。 我说，你会以“我父啊”称呼我， 不再转离而跟从我。
JER|3|20|以色列 家啊，你们向我行诡诈， 真像妻子行诡诈离开丈夫。 这是耶和华说的。
JER|3|21|有声音从光秃的高地传来， 就是 以色列 人哭泣恳求的声音， 因为他们走弯曲之道， 忘记耶和华－他们的上帝。
JER|3|22|“你们这背道的儿女啊，回来吧！ 我要医治你们背道的病。” “看哪，我们来到你这里， 因你是耶和华－我们的上帝。
JER|3|23|从小山来的真是枉然， 大山的喧嚷也是枉然 。 以色列 得救，诚然在乎耶和华－我们的上帝。
JER|3|24|“从我们幼年以来，那可耻之物 吞吃了我们祖先劳碌得来的，就是他们的羊群、牛群和他们的儿女。
JER|3|25|我们在羞耻中躺卧吧！愿惭愧将我们遮盖！因为从我们幼年以来，我们和我们的祖先都得罪了耶和华－我们的上帝，没有听从耶和华－我们上帝的话。”
JER|4|1|耶和华说：“ 以色列 啊， 你若回转，回转归向我， 若从我眼前除掉你可憎的偶像， 不再犹疑不定，
JER|4|2|凭诚实、公平、公义 指着永生的耶和华起誓； 列国就必因他蒙福， 也必因他夸耀。”
JER|4|3|耶和华对 犹大 人和 耶路撒冷 人如此说： “你们要为自己开垦荒地， 不要撒种在荆棘里。
JER|4|4|犹大 人和 耶路撒冷 的居民哪， 你们当自行割礼，归耶和华， 将你们心里的污秽 除掉； 免得我的愤怒因你们的恶行发作， 如火燃起， 甚至无人能熄灭！”
JER|4|5|你们要在 犹大 传扬， 在 耶路撒冷 宣告，说： “当在国中吹角，高声呼叫说： ‘你们当聚集！ 我们好进入坚固城！’
JER|4|6|应当向 锡安 竖立大旗。 逃吧，不要迟延， 因我必使灾祸与大毁灭从北方来到。
JER|4|7|有狮子从密林中上来， 是毁坏列国的。 它已动身出离本处， 要使你的地荒凉， 使你的城镇变为废墟，无人居住。
JER|4|8|因此，你们当腰束麻布，哭泣哀号， 因为耶和华的烈怒并未转离我们。”
JER|4|9|耶和华说：“到那时，君王和领袖的心要失丧，祭司都要惊奇，先知都要诧异。”
JER|4|10|我说：“哀哉！主耶和华啊，你真是大大欺哄这百姓和 耶路撒冷 ，说：‘你们必得平安。’其实刀剑已经抵住喉咙了！”
JER|4|11|那时，必有话对这百姓和 耶路撒冷 说：“来自旷野光秃高地的热风吹向我的百姓 ，不是为簸扬，也不是为扬净。
JER|4|12|又有一阵比这更大的风向我刮来；现在，我要向他们宣读我的判决。”
JER|4|13|看哪，他必如云涌上； 他的战车如旋风， 他的马比鹰更快。 我们有祸了！ 我们败落了！
JER|4|14|耶路撒冷 啊，你当洗去心中的恶， 使你可以得救。 恶念在你里面要存到几时呢？
JER|4|15|有声音从 但 传出， 有灾祸从 以法莲山 传来。
JER|4|16|你们当传给列国， 看哪，要向 耶路撒冷 报告： “有围攻的人从远方来到， 向 犹大 的城镇大声喊叫。
JER|4|17|他们包围 耶路撒冷 ， 好像看守田园的， 因为它背叛了我。 这是耶和华说的。
JER|4|18|你的作风和行为招惹这事； 这是你罪恶的结果， 实在是苦， 刺透了你的心！”
JER|4|19|我的肺腑啊，我的肺腑啊，我心疼痛！ 我的心在我里面烦躁不安。 我不能静默不言， 因我已听见角声和打仗的喊声。
JER|4|20|毁坏的信息不断传来， 因为全地荒废。 我的帐棚忽然毁坏， 我的幔子顷刻破裂。
JER|4|21|我看见大旗，听见角声， 要到几时呢？
JER|4|22|“我的百姓愚顽，不认识我； 他们是愚昧无知的儿女， 有智慧行恶，没有知识行善。”
JER|4|23|我观看地， 看哪，地是空虚混沌； 我观看天，天也无光。
JER|4|24|我观看大山，看哪，尽都震动， 小山也都摇来摇去。
JER|4|25|我观看，看哪，无人； 空中的飞鸟也都躲避。
JER|4|26|我观看，看哪，肥田变为荒地； 所有城镇在耶和华面前， 因他的烈怒都被拆毁。
JER|4|27|耶和华如此说：“全地必然荒凉， 我却不毁灭净尽。
JER|4|28|因此，地要悲哀， 天上也必黑暗； 因为我言已出，我意已定， 必不改变，也不由此转回。”
JER|4|29|各城的人因骑兵和弓箭手的响声就都逃跑， 进入密林，爬上磐石； 城镇都被抛弃， 无人住在其中。
JER|4|30|你这被毁灭的啊， 你要做什么呢？ 你穿上朱红衣服， 佩戴黄金饰物， 用眼影修饰眼睛， 徒然美化你自己。 恋慕你的却藐视你， 寻索你的性命。
JER|4|31|我听见仿佛妇人临产的声音， 好像生头胎疼痛的声音， 原来是 锡安 的声音； 她喘着气，伸开手： “我有祸了！ 在杀人者跟前，我的心灵发昏。”
JER|5|1|你们要走遍 耶路撒冷 的街市， 在广场寻找， 看是否有人行公平、求诚实； 若有，我就赦免这城。
JER|5|2|虽然他们说“我对永生的耶和华发誓”， 所起的誓实在是假的。
JER|5|3|耶和华啊，你的眼目不是在寻找诚实吗？ 你击打他们，他们却不伤恸； 你摧毁他们，他们仍不领受管教。 他们使脸刚硬过于磐石， 不肯回头。
JER|5|4|我说：“这些人实在是贫寒的， 他们是愚昧的， 因为不知道耶和华的作为， 也不知道他们上帝的法则。
JER|5|5|我要去见尊贵的人，向他们说话， 他们应该知道耶和华的作为， 知道他们上帝的法则。” 然而，这些人却齐心将轭折断， 挣开绳索。
JER|5|6|因此，林中的狮子必害死他们， 野地的狼必灭绝他们， 豹子在城外窥伺。 凡出城的必被撕碎， 因为他们的罪过极多， 背道的事也增加。
JER|5|7|我怎能赦免你呢？ 你的儿女离弃我， 又指着那不是上帝的起誓。 我使他们饱足， 他们就行奸淫， 居住 在娼妓家里。
JER|5|8|他们如喂饱的马，精力旺盛， 各向邻舍的妻子吹哨。
JER|5|9|我岂不因这些事施行惩罚吗？ 像这样的国家，我岂能不报复呢？ 这是耶和华说的。
JER|5|10|你们要上去毁坏它的葡萄园， 但不可毁坏净尽， 只可除掉其枝子， 因为不属耶和华。
JER|5|11|以色列 家和 犹大 家向我大行诡诈。 这是耶和华说的。
JER|5|12|关乎耶和华他们说了虚谎的话： “他不会的， 灾祸必不临到我们， 我们也不会遇见刀剑和饥荒。
JER|5|13|先知不过是一阵风， 道也不在他们里面； 这灾祸必临到他们身上。”
JER|5|14|所以耶和华－万军之上帝如此说： “因为他们说这话， 看哪，我必使我的话在你口中为火， 使这百姓为柴， 火便将他们烧灭。
JER|5|15|以色列 家啊， 看哪，我必使一国从远方来攻击你， 是强盛的国， 是古老的国； 他们的言语你不知道， 所说的话你不明白。 这是耶和华说的。
JER|5|16|他们的箭袋有如敞开的坟墓， 他们全都是勇士。
JER|5|17|他们必吃尽你的庄稼和粮食， 是你儿女该吃的 ； 必吃尽你的牛羊， 吃尽你的葡萄和无花果； 又必用刀剑毁坏你所倚靠的坚固城。
JER|5|18|“就是在那些日子，我也不会将你们毁灭净尽。这是耶和华说的。
JER|5|19|百姓若说：‘耶和华－我们的上帝为什么向我们行这一切事呢？’你就对他们说：‘你们怎样离弃我，在你们的地上事奉外邦神明，也必照样在不属你们的地上事奉外族人。’”
JER|5|20|当在 雅各 家传扬， 在 犹大 宣告，说：
JER|5|21|“愚昧无知的百姓啊， 你们有眼不看， 有耳不听， 现在当听这话。
JER|5|22|你们难道不惧怕我吗？ 在我面前还不战兢吗？ 这是耶和华说的。 我以沙为海的界限， 作永远的条例，使它不得越过。 波浪汹涌，却不能胜过； 怒涛澎湃，仍无法越过。
JER|5|23|但这百姓有背叛忤逆的心， 他们转离而去。
JER|5|24|他们心里并不说： ‘我们应当敬畏耶和华－我们的上帝； 他按时赐雨，就是秋雨和春雨， 又为我们定收割的季节。’
JER|5|25|你们的罪孽使这些转离你们， 你们的罪恶使你们不能得福。
JER|5|26|在我百姓当中有恶人， 他们埋伏，好像捕鸟的人在窥探 ； 他们设罗网陷害人。
JER|5|27|笼子怎样装满雀鸟， 他们的屋里也照样充满诡诈； 他们因此得以强大富足。
JER|5|28|他们肥胖光润，作恶过甚， 不为人伸冤， 不为孤儿伸冤，使他们胜诉， 也不为贫穷人辩护。
JER|5|29|我岂不因这些事施行惩罚吗？ 像这样的国家，我岂能不报复呢？ 这是耶和华说的。
JER|5|30|“国中有令人惊骇、 恐怖的事发生，
JER|5|31|先知说假预言， 祭司把权柄抓在自己手上， 我的百姓也喜爱这样， 到了结局你们要怎么办呢？”
JER|6|1|便雅悯 人哪，当逃离 耶路撒冷 ， 在 提哥亚 吹号角， 在 伯．哈基琳 升信号， 因为有灾祸与大毁灭从北方逼近。
JER|6|2|那秀美娇嫩的 锡安 ， 我必剪除。
JER|6|3|牧人必引领羊群到它那里， 在它周围支搭帐棚， 各在自己的地方放牧。
JER|6|4|“你们要准备攻击它。 起来吧，我们要趁正午上去。” “哀哉！日已渐斜， 黄昏的影子拖长了。”
JER|6|5|“起来吧，我们要在夜间上去， 毁坏它的宫殿。”
JER|6|6|万军之耶和华如此说： “你们要砍伐树木， 建土堆攻打 耶路撒冷 ， 就是那该受罚的城 ， 其中尽是欺压。
JER|6|7|井怎样涌出水来， 这城也照样涌出恶来； 其中常听闻残暴毁灭的事， 病痛损伤也常在我面前。
JER|6|8|耶路撒冷 啊，当受管教， 免得我心与你生疏， 免得我使你荒凉， 成为无人居住之地。”
JER|6|9|万军之耶和华如此说： “他们洗劫 以色列 剩下的民， 如摘净葡萄一样； 现你的手如采收葡萄的人，在树枝上采了又采 。”
JER|6|10|现在我可以向谁说话，警告谁，使他们听呢？ 看哪，他们的耳朵未受割礼，不能听见。 看哪，他们以耶和华的话为羞辱， 不以为喜悦。
JER|6|11|因此我被耶和华的愤怒充满，难以忍受。 “你要把它倒在街上孩童 和成群的年轻人身上， 他们连夫带妻， 年长者与高龄的人都必被擒拿。
JER|6|12|他们的房屋、田地， 和妻子都要一起转归别人， 我要伸手攻击这地的居民。” 这是耶和华说的。
JER|6|13|“因为他们从最小的到最大的都贪图不义之财， 从先知到祭司全都行事虚假。
JER|6|14|他们轻忽地医治我百姓的损伤， 说：‘平安了！平安了！’ 其实没有平安。
JER|6|15|他们行可憎之事，应当羞愧； 然而他们却一点也不觉得羞愧， 也不知羞耻。 因此，他们必与仆倒的人一同仆倒， 我惩罚他们的时候， 他们必跌倒。” 这是耶和华说的。
JER|6|16|耶和华如此说： “你们当站在路边察看， 寻访古老的路， 哪里是完善的道路，就行走在其上； 这样，你们自己必找到安息。 他们却说：‘我们不走。’
JER|6|17|我为你们设立守望的人， 要留心听角声。 他们却说：‘我们不听。’
JER|6|18|因此，列国啊，当听！ 会众啊，要知道他们必遭遇的事。
JER|6|19|地啊，当听！ 看哪，我必使灾祸临到这百姓， 是他们计谋所结的果子； 因为他们不肯留心听我的话， 至于我的律法，他们也厌弃。
JER|6|20|从 示巴 来的乳香， 从远方出的香菖蒲， 奉来给我有何用呢？ 你们的燔祭不蒙悦纳； 你们的祭物，我也不喜悦。”
JER|6|21|所以耶和华如此说： “看哪，我要将绊脚石放在这百姓面前； 父亲和儿子要一同跌在其上， 邻舍与朋友也都灭亡。”
JER|6|22|耶和华如此说： “看哪，有一民族从北方而来； 有一大国被激起，从地极来到。
JER|6|23|他们拿弓和枪， 性情残忍，不施怜悯； 他们的声音如海浪澎湃。 锡安 哪， 他们都骑马， 如上战场的人摆阵攻击你。”
JER|6|24|我们听见这样的风声，手就发软； 痛苦将我们抓住， 疼痛仿佛临产的妇人。
JER|6|25|你们不要出到田野去， 也不要行走在路上， 因四围有仇敌的刀剑和惊吓。
JER|6|26|我的百姓 啊，应当腰束麻布，滚在灰中。 要悲伤，如丧独子般痛痛哭号， 因为灭命的忽然临到我们。
JER|6|27|我使你作我百姓的测试者 和考验者 ， 使你知道并考验他们的行为。
JER|6|28|他们极其悖逆， 到处毁谤人， 他们是铜是铁， 全都败坏了。
JER|6|29|风箱吹火，铅被烧毁， 炼而又炼，终是徒然， 因为恶劣的还未除掉。
JER|6|30|人必称他们为被抛弃的银子， 因为耶和华已经抛弃了他们。
JER|7|1|耶和华的话临到 耶利米 ，说：
JER|7|2|“你当站在耶和华殿的门口，在那里宣讲这话说：所有从这些门进来敬拜耶和华的 犹大 人哪，当听耶和华的话。
JER|7|3|万军之耶和华－ 以色列 的上帝如此说：你们要改正你们的所作所为，我就使你们仍然居住这地 。
JER|7|4|不要倚靠虚谎的话，说：‘这是耶和华的殿，是耶和华的殿，是耶和华的殿！’
JER|7|5|“你们若实在改正你们的所作所为，彼此诚然施行公平，
JER|7|6|不欺压寄居的和孤儿寡妇，不在这地方流无辜人的血，也不随从别神陷害自己，
JER|7|7|我就使你们仍然居住这地 ，就是我从古时所赐给你们祖先的地，从永远到永远。
JER|7|8|“看哪，你们倚靠虚谎无益的话语。
JER|7|9|你们岂可偷盗，杀害，奸淫，起假誓，向 巴力 烧香，随从素不认识的别神，
JER|7|10|又来到这称为我名下的殿，在我面前敬拜，说‘我们平安无事’，为了要行这一切可憎的事呢？
JER|7|11|这称为我名下的殿在你们眼中岂可看为贼窝呢？看哪，我真的都看见了。这是耶和华说的。
JER|7|12|你们到我的地方 示罗 去，就是我先前在那里立为我名的居所，察看我因这百姓 以色列 的罪恶向那地方所行的事。
JER|7|13|现在，因你们行了这一切的事，我一再警戒你们，你们却不听从；我呼唤你们，你们也不回应。这是耶和华说的。
JER|7|14|所以我要向这称为我名下、你们所倚靠的殿，与我所赐给你们和你们祖先的地这样行，正如我从前向 示罗 所行的。
JER|7|15|我必将你们从我眼前赶出，正如赶出你们的众弟兄，就是所有 以法莲 的后裔。”
JER|7|16|“所以，你不要为这百姓祈祷；不要为他们呼求祷告，也不要为他们向我祈求，因我不听你。
JER|7|17|他们在 犹大 城镇和 耶路撒冷 街上所做的，你难道没有看见吗？
JER|7|18|孩子捡柴，父亲烧火，妇女揉面做饼，献给天后，又向别神献浇酒祭，惹我发怒。
JER|7|19|他们岂是惹我发怒呢？不是自己惹祸，以致脸上惭愧吗？这是耶和华说的。
JER|7|20|所以主耶和华如此说：看哪，我必将我的怒气和愤怒倾倒在这地方的人和牲畜身上、田野的树木和地里的出产上，它必燃烧，不会熄灭。”
JER|7|21|万军之耶和华－ 以色列 的上帝如此说：“你们要将燔祭加在你们的祭物上，又要吃肉；
JER|7|22|因为我将你们祖先从 埃及 地领出来的那日，燔祭和祭物的事我并没有提说，也没有吩咐他们。
JER|7|23|我只吩咐他们这一件事说：‘你们当听从我的话，我就作你们的上帝，你们也作我的子民。你们行走我所吩咐的一切道路，就可以得福。’
JER|7|24|他们却不听从，也不侧耳而听，竟随从自己的计谋和顽梗的恶心去行，不进反退。
JER|7|25|自从你们祖先出 埃及 地的那日，直到今日，我每日一再差遣我的仆人众先知到你们那里去。
JER|7|26|你们却不听我，不侧耳而听，竟硬着颈项行恶，比你们的祖先更甚。
JER|7|27|“你要将这一切的话告诉他们，他们却不听你；呼唤他们，他们却不回应。
JER|7|28|你要对他们说：‘这就是不听从耶和华－他们上帝的话、不领受训诲的国民；诚信已从他们口中消失殆尽了。
JER|7|29|耶路撒冷 啊，要剪头发，扔掉它， 在光秃的高地唱哀歌， 因为耶和华弃绝、离弃了惹他发怒的世代。’”
JER|7|30|“ 犹大 人行我眼中看为恶的事，将可憎之偶像立在称为我名下的殿里，玷污这殿。这是耶和华说的。
JER|7|31|他们在 欣嫩子谷 建造 陀斐特 的丘坛，要在火中焚烧自己的儿女。这并不是我所吩咐的，我心里也从来没有想过。
JER|7|32|因此，看哪，日子将到，这地方不再称为 陀斐特 和 欣嫩子谷 ，反倒称为 杀戮谷 。他们要在 陀斐特 埋葬尸首，甚至无处可葬。这是耶和华说的。
JER|7|33|并且这百姓的尸首要给空中的飞鸟和地上的走兽作食物，无人吓走它们。
JER|7|34|那时，我必止息 犹大 城镇和 耶路撒冷 街上欢喜和快乐的声音、新郎和新娘的声音，因为这地必然荒芜。”
JER|8|1|耶和华说：“那时，人必将 犹大 诸王和领袖的骸骨、祭司和先知的骸骨，以及 耶路撒冷 居民的骸骨，都从坟墓中取出来，
JER|8|2|散布在太阳、月亮和天上众星之下，就是他们从前所喜爱、所事奉、所随从、所求问、所敬拜的。这些骸骨不被收殓，不被埋葬，必在地面上成为粪土。
JER|8|3|这邪恶家族所幸存的余民，就是在我赶他们到的各处所剩下的 ，全都宁可选死不选活。这是万军之耶和华说的。”
JER|8|4|“你要对他们说，耶和华如此说： 人跌倒，不再起来吗？ 人转去，不再转回来吗？
JER|8|5|这 耶路撒冷 的百姓为何永久背道呢？ 他们抓住诡诈，不肯回头。
JER|8|6|我留心听，听见他们说不诚实的话。 无人懊悔自己的恶行，说： ‘我做的是什么呢？’ 他们全都转奔己路， 如马直闯战场。
JER|8|7|空中的鹳鸟知道自己的季节， 斑鸠、燕子与白鹤也守候当来的时令； 我的百姓却不知道耶和华的法则。
JER|8|8|“你们怎么说：‘我们有智慧， 耶和华的律法在我们这里’？ 看哪，其实文士的假笔舞弄虚假。
JER|8|9|智慧人惭愧，惊惶，被擒拿； 看哪，他们背弃耶和华的话， 还会有什么智慧呢？
JER|8|10|因此，我必将他们的妻子给别人， 将他们的田地给别人为业； 因为他们从最小的到最大的都贪图不义之财， 从先知到祭司全都行事虚假。
JER|8|11|他们轻忽地医治我百姓的损伤，说： ‘平安了！平安了！’ 其实没有平安。
JER|8|12|他们行可憎之事，应当羞愧； 然而他们却一点也不觉得羞愧， 又不知羞耻。 因此，他们必与仆倒的人一样仆倒； 我惩罚他们的时候， 他们必跌倒。 这是耶和华说的。
JER|8|13|我必使他们全然灭绝； 葡萄树上必没有葡萄 ， 无花果树上没有果子， 叶子也必枯干。 我所赐给他们的， 必离他们而去。 这是耶和华说的。”
JER|8|14|我们为何静坐不动呢？ 我们当聚集，进入坚固城， 在那里静默不言； 因为耶和华－我们的上帝使我们静默不言， 又将苦水给我们喝， 都因我们得罪了耶和华。
JER|8|15|我们指望平安， 却得不着福气； 指望痊愈的时刻， 看哪，受了惊惶。
JER|8|16|“从 但 那里传来敌人的马喷气的声音， 壮马发出嘶声， 全地就都震动； 因为他们来吞灭这地和其上所有的， 吞灭这城与其中的居民。
JER|8|17|看哪，我必派蛇进到你们中间， 就是法术无法驱除的毒蛇， 它们必咬你们。 这是耶和华说的。”
JER|8|18|忧愁时我寻找安慰 ， 我心在我里面发昏。
JER|8|19|听啊，是我百姓呼救的声音从远地传来： “耶和华不是在 锡安 吗？ 锡安 的王不是在其中吗？” “他们为什么以自己雕刻的偶像 和外邦虚无的神明 惹我发怒呢？”
JER|8|20|“秋收已过，夏季已完， 我们还未得救！”
JER|8|21|因我百姓的损伤， 我也受了损伤。 我哀恸，惊惶将我抓住。
JER|8|22|在 基列 岂没有乳香呢？ 在那里岂没有医生呢？ 我百姓 为何得不着医治呢？
JER|9|1|但愿我的头为水， 我的眼为泪水的泉源， 我好为我百姓 中被杀的人昼夜哭泣。
JER|9|2|惟愿在旷野有旅客的客栈， 我好离开我的百姓而去； 因他们全都行奸淫， 是行诡诈的一党。
JER|9|3|他们弯起舌头像弓， 为要说谎话； 他们在国中增长势力， 不是为诚信。 他们恶上加恶， 并不认识我。 这是耶和华说的。
JER|9|4|你们各人当谨防邻舍， 不可信赖弟兄； 因为弟兄尽行欺骗， 邻舍也都往来毁谤人。
JER|9|5|他们互相欺骗， 不说真话， 训练自己的舌头说谎， 竭尽所能地作恶。
JER|9|6|你居住在诡诈的人中； 他们因行诡诈 ，不愿意认识我。 这是耶和华说的。
JER|9|7|所以万军之耶和华如此说： “看哪，我要熬炼他们，考验他们； 不然，为了我的百姓 ，我该如何行呢？
JER|9|8|他们的舌头是毒箭，说话诡诈， 跟邻舍口说平安， 心却谋害他。
JER|9|9|我岂不因这些事向他们施行惩罚吗？ 像这样的国家，我岂能不报复呢？ 这是耶和华说的。”
JER|9|10|我要为山岭哭泣悲哀， 为旷野的草场扬声哀号； 因为都已枯焦，甚至无人经过。 牲畜的鸣叫听不见， 空中的飞鸟和地上的走兽也都逃离。
JER|9|11|我必使 耶路撒冷 成为废墟，为野狗的住处， 也必使 犹大 的城镇荒废，无人居住。
JER|9|12|谁是智慧人，可以明白这事？耶和华的口可向谁述说，使他传讲呢？这地为何毁灭，枯焦如旷野，无人经过呢？
JER|9|13|耶和华说：“因为这百姓离弃我在他们面前所设立的律法，不听从我的话，不肯遵行，
JER|9|14|反随从自己顽梗的心行事，照他们祖先所教训的随从诸 巴力 。”
JER|9|15|所以万军之耶和华－ 以色列 的上帝如此说：“看哪，我必将茵蔯给这百姓吃，又用苦水给他们喝。
JER|9|16|我要把他们分散在他们和他们祖宗所不认识的列国；我也要使刀剑追杀他们，直到将他们灭尽。”
JER|9|17|万军之耶和华如此说： “你们要考虑， 将唱哀歌的妇女召来， 差人召善哭的妇女前来，
JER|9|18|叫她们速速为我们举哀， 使我们泪眼汪汪， 使我们的眼皮涌出泪水。
JER|9|19|因为有哀声从 锡安 传来： ‘我们竟然败落！ 我们何等惭愧！ 我们撇下土地， 人拆毁了我们的房屋。’”
JER|9|20|妇女们哪，当听耶和华的话， 领受他口中的言语； 当教导你们的女儿举哀， 各人教导女伴唱哀歌。
JER|9|21|因为死亡从窗户进来， 进入我们的宫殿， 从外边剪除孩童， 从街上剪除少年。
JER|9|22|你当说，耶和华如此说： 人的尸首必倒在田野像粪土， 又像收割的人身后遗落的禾稼， 无人拾取。
JER|9|23|耶和华如此说：“智慧人不要因他的智慧夸口，勇士不要因他的力气夸口，财主也不要因他的财富夸口；
JER|9|24|夸口的却要夸自己有聪明，认识我是耶和华，知道我喜悦在世上施行慈爱、公平和公义。这是耶和华说的。
JER|9|25|“看哪，日子将到，这是耶和华说的，我要惩罚只在肉身受割礼的人，
JER|9|26|就是 埃及 、 犹大 、 以东 、 亚扪 人、 摩押 人，和住旷野所有剃鬓发的人；因为列国都未受割礼， 以色列 全家心中也未受割礼。”
JER|10|1|以色列 家啊，要听耶和华对你们所说的话，
JER|10|2|耶和华如此说： “不要效法列国的行为， 任凭列国因天象惊惶， 你们不要惊惶。
JER|10|3|万民的习俗是虚空的； 偶像 不过是从树林中砍来的木头， 是匠人用斧头做成的手工。
JER|10|4|人用金银妆饰它， 用钉子和锤子钉稳， 使它不动摇。
JER|10|5|偶像好像瓜田里的稻草人， 不能说话，不能行走， 必须有人抬着。 不要怕它们， 因它们不能降祸， 也无力降福。”
JER|10|6|耶和华啊，没有谁能与你相比！ 你本为大，你的名也大有能力。
JER|10|7|万国的王啊，谁不敬畏你？ 敬畏你本是合宜的； 列国所有的智慧人中， 在他们一切的国度里， 都没有能与你相比的。
JER|10|8|他们如同畜牲，尽都愚昧。 偶像的训诲算什么呢？ 偶像不过是木头，
JER|10|9|锤炼的银片是从 他施 来的， 金子则从 乌法 而来， 都是匠人和银匠的手工； 又有蓝色和紫色的衣服， 全都是巧匠的作品。
JER|10|10|惟耶和华是真上帝， 是活的上帝，是永远的王。 他一发怒，大地震动； 他一恼恨，列国担当不起。
JER|10|11|你们要对他们这样说：“那些不是创造天地的神明，必从地上、从天下被除灭！”
JER|10|12|耶和华以能力创造大地， 以智慧建立世界， 以聪明铺张穹苍。
JER|10|13|他一出声，天上就有众水澎湃； 他使云雾从地极上腾， 造电随雨而闪， 从仓库中吹出风来。
JER|10|14|人人都如同畜牲，毫无知识； 银匠都因偶像羞愧， 他所铸的偶像本是虚假， 它们里面并无气息。
JER|10|15|偶像都是虚无的， 是迷惑人的作品， 到受罚的时刻必被除灭。
JER|10|16|雅各 所得的福分不是这样， 因主 是那创造万有的， 以色列 是他产业的支派， 万军之耶和华是他的名。
JER|10|17|受围困的居民哪，当收拾你的行囊， 离开这地。
JER|10|18|因为耶和华如此说： “看哪，这一次，我必将此地的居民抛出去， 又必加害他们， 使他们觉悟 。”
JER|10|19|祸哉！我受损伤， 我的伤痕极其重大。 我却说：“这真的是我必须忍受的痛苦。”
JER|10|20|我的帐棚毁坏， 我的绳索折断， 我的儿女都离我而去，不在了。 再无人来支搭我的帐棚，挂起我的幔子。
JER|10|21|因为牧人如同畜牲， 没有寻求耶和华， 所以不得顺利； 他们的羊群也都分散了。
JER|10|22|有风声！看哪，来了！ 有大扰乱从北方而来， 要使 犹大 的城镇变为废墟， 成为野狗的住处。
JER|10|23|耶和华啊，我知道人的道路不由自己， 行路的人也不能定自己的脚步。
JER|10|24|耶和华啊，求你按公平管教我， 不要在你的怒中惩治我， 免得你使我归于无有。
JER|10|25|求你将愤怒倾倒在不认识你的列国中， 倾倒在不求告你名的各族上； 因为他们吞了 雅各 ，不但吞吃，而且灭绝， 使他的住处变为荒凉。
JER|11|1|耶和华的话临到 耶利米 ，说：
JER|11|2|“当听这约的话，告诉 犹大 人和 耶路撒冷 的居民，
JER|11|3|对他们说，耶和华－ 以色列 的上帝如此说：‘不听从这约之话的人必受诅咒。
JER|11|4|这约是我将你们祖先从 埃及 地领出来，脱离铁炉的那日所吩咐他们的，说：你们要听从我的话，照我所吩咐的一切去做。这样，你们作我的子民，我也作你们的上帝，
JER|11|5|我好坚定我向你们列祖所起的誓，赏赐他们流奶与蜜之地，正如今日一样。’”我就回应说：“耶和华啊，阿们！”
JER|11|6|耶和华对我说：“你要在 犹大 城镇和 耶路撒冷 街市宣告这一切话，说：‘当听从遵行这约的话，
JER|11|7|因为我将你们祖先从 埃及 地领出来的那日，直到今日，都一再切切告诫他们说：当听从我的话。
JER|11|8|他们却不听从，也不侧耳而听，竟随从自己顽梗的恶心去行。我就使这约中一切诅咒的话临到他们身上；这约是我吩咐他们遵行的，他们却不遵行。’”
JER|11|9|耶和华对我说：“在 犹大 人和 耶路撒冷 居民中有同谋背叛的事。
JER|11|10|他们转去效法他们祖先的恶行，不肯听我的话，竟随从别神，事奉它们。 以色列 家和 犹大 家违背了我与他们列祖所立的约。
JER|11|11|所以耶和华如此说：看哪，我必使灾祸临到他们，是他们不能逃脱的。他们向我哀求，我却不听。
JER|11|12|那时， 犹大 城镇的人和 耶路撒冷 的居民要哀求他们烧香所供奉的神明；只是遭难的时候，这些神明一点也不能拯救他们。
JER|11|13|犹大 啊，你神明的数目与你城镇的数目相等；你所筑可耻的坛，就是向 巴力 烧香的坛 ，也与 耶路撒冷 街道的数目相等。
JER|11|14|“所以你不要为这百姓祈祷，也不要为他们呼求祷告，因为他们遭难向我哀求的时候，我必不应允。
JER|11|15|我所亲爱的既多设恶谋，还能在我殿中做什么呢？你因作恶就喜乐，圣肉要离开你。
JER|11|16|从前耶和华给你起名叫青橄榄树，又华美又结好果子；如今他用一声巨响点火在其上，枝子就折断了。
JER|11|17|“原来栽培你的万军之耶和华已经说要降祸给你，是因 以色列 家和 犹大 家行恶。他们向 巴力 烧香，惹我发怒，是自作自受。”
JER|11|18|耶和华指示我，我才知道； 你将他们所做的给我指明。
JER|11|19|我像柔顺的羔羊被牵去宰杀， 并不知道他们设计谋害我： “我们把树连果子都灭了吧！ 把他从活人之地剪除， 使他的名不再被记得。”
JER|11|20|按公义判断、察验人肺腑心肠的万军之耶和华啊， 求你使我得见你在他们身上报仇， 因我已将我的案件向你禀明了。
JER|11|21|所以，耶和华论到寻索你命的 亚拿突 人如此说：“他们说：你不要奉耶和华的名说预言，免得你死在我们手中。
JER|11|22|所以万军之耶和华如此说：看哪，我必惩罚他们；他们的壮丁必被刀剑杀死，他们的儿女必因饥荒而死，
JER|11|23|他们当中必无任何幸存者；因为在他们受罚之年，我必使灾祸临到 亚拿突 人。”
JER|12|1|耶和华啊，我与你争辩的时候， 你总是显为义； 但有一件，我还要与你理论： 恶人的道路为何亨通呢？ 大行诡诈的为何得安逸呢？
JER|12|2|你栽培了他们， 他们也扎了根， 长大，而且结果。 他们的口与你相近， 心却与你远离。
JER|12|3|耶和华啊，你认识我，看见我， 你察验我向你的心如何。 求你将他们拉出来， 如将宰的羊， 为杀戮的日子分别出来。
JER|12|4|这地悲哀， 一切田野的青草枯干要到几时呢？ 因其上居民的恶行， 牲畜和飞鸟都灭绝了。 因为他们说：“他看不见 我们的结局 。”
JER|12|5|“你与步行的人同跑， 尚且觉得累， 怎能与马赛跑呢？ 你在安全之地尚且会跌倒 ， 在 约旦河 边的丛林要怎么办呢？
JER|12|6|因为连你兄弟和你父家都以诡诈待你， 甚至在你后边大声喊叫。 虽然他们向你说好话， 你也不要相信他们。”
JER|12|7|我离弃了我的殿宇， 撇弃了我的产业， 将我心里所亲爱的交在她 仇敌手中。
JER|12|8|我的产业向我如林中的狮子， 出声攻击我， 因此我恨恶她。
JER|12|9|我的产业向我如斑点的鸷鸟， 有鸷鸟在四围攻击她。 你们去聚集田野的百兽， 叫它们来吞吃吧！
JER|12|10|许多牧人毁坏我的葡萄园， 践踏我的地产， 使我美好的地产变为荒凉的旷野。
JER|12|11|他们使地荒凉； 地既荒凉，就向我哀哭。 全地荒凉，却无人在意。
JER|12|12|灭命的来到旷野中一切光秃的高地； 耶和华的刀从地这边直到地那边，尽行杀灭， 凡血肉之躯都不得平安。
JER|12|13|他们种的是麦子， 收的却是荆棘； 辛辛苦苦却无收获。 因耶和华的烈怒， 你们必为自己的收成感到羞愧。
JER|12|14|耶和华如此说：“看哪，我要将所有的恶邻拔出本地，他们曾占据了我赐给 以色列 百姓所承受的产业；我也要将 犹大 家从他们中间拔出来。
JER|12|15|我拔出他们以后，必回转过来怜悯他们，使他们归回，各归本业，各归故土。
JER|12|16|他们若殷勤学习我百姓的道，指着我的名起誓：‘我指着永生的耶和华起誓’，正如他们从前教我百姓指着 巴力 起誓，他们必在我百姓中得以建立。
JER|12|17|他们若是不听，我必拔出那国，不但拔出，还要毁灭。这是耶和华说的。”
JER|13|1|耶和华对我如此说：“你去买一条麻布带子，束在你腰上，不可把它泡在水里。”
JER|13|2|我就照耶和华的话，买了一条带子，束在我的腰上。
JER|13|3|耶和华的话第二次临到我，说：
JER|13|4|“要拿你所买、在你腰上的带子，起来往 幼发拉底河 去，把腰带藏在那里的磐石穴中。”
JER|13|5|我就去，照着耶和华命令我的，把腰带藏在 幼发拉底河 边。
JER|13|6|过了多日，耶和华对我说：“你起来往 幼发拉底河 去，把我命令你藏在那里的腰带取出来。”
JER|13|7|我就往 幼发拉底河 去，把那腰带从我所藏的地方挖出来。看哪，腰带已经破烂，毫无用处了。
JER|13|8|耶和华的话临到我，说：
JER|13|9|“耶和华如此说：我要照样败坏 犹大 的骄傲和 耶路撒冷 的狂傲。
JER|13|10|这恶民不肯听我的话，按自己顽梗的心而行，随从别神，事奉敬拜它们；这恶民必像这腰带，毫无用处。
JER|13|11|腰带怎样紧贴人的腰，照样，我也曾使 以色列 全家和 犹大 全家紧贴着我，归我为子民，使我得名声，得颂赞，得荣耀；他们却不肯听从。这是耶和华说的。”
JER|13|12|“所以你要对他们说：‘耶和华－ 以色列 的上帝如此说：各坛都要装满酒。’他们必对你说：‘我们岂不知道各坛都要装满酒吗？’
JER|13|13|你就对他们说：‘耶和华如此说：看哪，我必使这地所有的居民，就是坐 大卫 宝座的君王、祭司和先知，并 耶路撒冷 所有的居民，都酩酊大醉。
JER|13|14|我要使他们彼此冲突，连父与子也互相冲突；我必不可怜，不顾惜，不怜悯，以致将他们灭绝。这是耶和华说的。’”
JER|13|15|你们当听，当侧耳而听； 不可骄傲，因为耶和华已经吩咐了。
JER|13|16|当耶和华－你们的上帝 尚未使黑暗来临， 在昏暗的山上 你们的脚未绊跌以前， 要将荣耀归给他。 你们盼望光明， 他却使光明变为死荫， 成为幽暗。
JER|13|17|你们若不听这话， 我的心必因你们的骄傲暗自哭泣； 我的眼必痛哭流泪， 因为耶和华的羊群被掳去了。
JER|13|18|你要对君王和太后说： “你们当自卑，坐下； 因你们的王冠， 就是你们华美的冠冕已经掉落了 。”
JER|13|19|尼革夫 的城镇都被关闭， 无人打开； 犹大 全被掳掠， 掳掠净尽。
JER|13|20|你们要举目观看从北方来的人。 先前赐给你的羊群， 就是你所引以为荣的羊， 现今在哪里呢？
JER|13|21|耶和华立你自己所教导的盟友， 立他们为头来辖制你， 你还有什么话可说呢？ 痛苦岂不将你抓住像临产的妇人吗？
JER|13|22|你若心里说：“这一切的事为何临到我呢？” 是因你罪孽甚多。 你的下摆揭起， 你的脚跟受伤。
JER|13|23|古实 人岂能改变皮肤呢？ 豹岂能改变斑点呢？ 若能，你们这善于行恶的便能行善了。
JER|13|24|我必吹散他们， 如碎秸随旷野的风飘动。
JER|13|25|这是你所当得的， 是我量给你的报应 ； 因为你忘记了我， 倚靠虚假 。 这是耶和华说的。
JER|13|26|我要揭起你的下摆， 蒙在你脸上， 显露你的羞耻。
JER|13|27|你在田野的山上行奸淫， 发嘶声，谋淫乱， 这些可憎之事我都看见了。 耶路撒冷 啊，你有祸了！ 你不肯洁净 还要等到几时呢？
JER|14|1|耶和华的话临到 耶利米 ，论到旱灾的事：
JER|14|2|“ 犹大 悲哀，城门衰败； 众人坐在地上哀恸， 耶路撒冷 的哀声上达。
JER|14|3|他们的贵族打发童仆去打水； 他们来到水池， 找不到水，就拿着空器皿， 蒙羞惭愧，抱头而回。
JER|14|4|因为无雨降在地上，土地就干裂， 农夫为此蒙羞抱头。
JER|14|5|田野的母鹿因为无草 也撇弃才生的小鹿。
JER|14|6|野驴站在光秃的高地喘气，好像野狗； 它们的眼目因无草而失明。”
JER|14|7|耶和华啊，虽然我们的罪孽控告我们， 求你为你名的缘故行动吧！ 我们本是多次背道，得罪了你。
JER|14|8|以色列 所盼望，在患难时作他救主的啊， 你在这地为何像寄居的， 又如旅行的只住一夜呢？
JER|14|9|你为何像受惊吓的人， 像不能救人的勇士呢？ 耶和华啊，你在我们中间， 我们是称为你名下的人， 求你不要离开我们。
JER|14|10|耶和华论到这百姓如此说： “这百姓喜爱游荡， 不约束自己的脚步， 所以耶和华不悦纳他们。 现今他要记起他们的罪孽， 惩罚他们的罪恶。”
JER|14|11|耶和华又对我说：“不要为这百姓求福。
JER|14|12|他们禁食的时候，我不听他们的呼求；他们献燔祭和素祭，我也不悦纳。我却要用刀剑、饥荒、瘟疫灭绝他们。”
JER|14|13|我就说：“唉！主耶和华，看哪，那些先知常对他们说：‘你们必不见刀剑，也不遭饥荒；耶和华要在这地方赏赐你们真正的平安。’”
JER|14|14|耶和华对我说：“那些先知托我的名说假预言，我并未差遣他们，没有吩咐他们，也没有对他们说话；他们向你们预言的是虚假的异象、占卜、虚无，以及心中的诡诈。
JER|14|15|所以耶和华如此说：‘论到托我名说预言的那些先知，我并未差遣他们；他们说这地不会有刀剑、饥荒，其实那些先知自己必被刀剑、饥荒灭绝。
JER|14|16|听他们说预言的百姓必因饥荒、刀剑被扔在 耶路撒冷 的街道上，无人埋葬。他们连妻子带儿女，都是如此。我必将他们的恶倒在他们身上。’”
JER|14|17|你要向他们说这些话： 愿我眼泪汪汪， 昼夜不息， 因为少女─我百姓 受了重大的打击， 伤口极其严重。
JER|14|18|我若出到田间， 看哪，有被刀杀的； 我若进入城内， 看哪，有因饥荒患病的； 先知和祭司也在各地往来经商， 不知如何是好。
JER|14|19|你全然弃绝 犹大 吗？ 你的心厌恶 锡安 吗？ 你为何击打我们，使我们无法得医治呢？ 我们指望平安，却得不着福气； 指望痊愈，看哪，受了惊惶。
JER|14|20|耶和华啊，我们承认自己的罪恶 和我们祖先的罪孽， 因我们得罪了你。
JER|14|21|求你为你名的缘故， 不厌恶，不轻视你荣耀的宝座。 求你记念， 不要违背你与我们所立的约。
JER|14|22|外邦虚无的神明 中有能降雨的吗？ 天能自降甘霖吗？ 耶和华－我们的上帝啊，不是你吗？ 我们要等候你， 因为这一切都是你所造的。
JER|15|1|耶和华对我说：“虽有 摩西 和 撒母耳 站在我面前，我的心也不顾惜这百姓。你把他们从我眼前赶出，叫他们出去吧！
JER|15|2|他们若问你说：‘我们往哪里去呢？’你就告诉他们，耶和华如此说： ‘定为死亡的，必致死亡； 定为刀杀的，必被刀杀； 定为饥荒的，必遭饥荒； 定为掳掠的，必被掳掠。’”
JER|15|3|“我命定四样灾害临到他们，就是刀剑杀戮、群狗拖拉、空中的飞鸟和地上的走兽吞吃毁灭。这是耶和华说的。
JER|15|4|我必使地上万国因他们而惊骇，都因 希西家 的儿子 犹大 王 玛拿西 在 耶路撒冷 所做的事。”
JER|15|5|耶路撒冷 啊，有谁同情你呢？ 有谁为你悲伤呢？ 有谁转身问你安呢？
JER|15|6|你弃绝了我， 转身退后； 因此我伸手攻击你，毁灭你， 我已怜悯到厌烦了。 这是耶和华说的。
JER|15|7|我在境内各关口 用簸箕筛我的百姓， 使他们丧掉儿女， 又毁灭他们， 他们仍不转离所行的道。
JER|15|8|他们的寡妇在我面前比海沙更多； 我使灭命者在正午来到， 攻击年轻人的母亲， 使痛苦惊吓忽然临到她身上。
JER|15|9|生过七个孩子的妇人衰弱； 尚在白昼，太阳忽然落下， 她就抱愧蒙羞。 我必当着敌人的面， 将他们当中的幸存者交给刀剑。 这是耶和华说的。
JER|15|10|我的母亲哪，我有祸了！因你生我作全地争相指控的人。我素来没有借贷给人，人也没有借贷给我，人人却都咒骂我。
JER|15|11|耶和华说：“我必定释放 你，使你得福气。灾祸苦难来临时，我必使仇敌央求你。
JER|15|12|人岂能将铜与铁，就是北方的铁折断呢？
JER|15|13|“我必因你在四境之内所犯的一切罪，将你的货物财宝当掠物，白白地交出来 。
JER|15|14|我要使你的仇敌过去，到你所不认识的地方 ，因为你们要被我怒中所起的火焚烧。”
JER|15|15|耶和华啊，你是知道的； 求你记念我，眷顾我， 向迫害我的人为我报仇； 不要把我取去，因你不轻易发怒， 要知道我为你的缘故受了凌辱。
JER|15|16|耶和华－万军之上帝啊， 我得着你的话就把它们吃了， 你的话是我心中的欢喜快乐； 因我是称为你名下的人。
JER|15|17|我并未坐在享乐人的会中欢乐； 因你的手，我就独自静坐， 你使我满心愤慨。
JER|15|18|我的痛苦为何长久不止呢？ 我的伤痕为何无法可医，不能痊愈呢？ 难道你以诡诈待我，像流干的河道吗？
JER|15|19|所以耶和华如此说：“你若回转， 我就使你归回， 站在我面前。 你若能将宝物和无用之物分别出来， 你就可以当作我的口。 他们必归向你， 你却不可归向他们。
JER|15|20|我必使你向这百姓成为坚固的铜墙。 他们必攻击你，却不能胜过你； 因我与你同在，要拯救你，搭救你。 这是耶和华说的。
JER|15|21|我必搭救你脱离恶人的手， 救赎你脱离残暴之人的手。”
JER|16|1|耶和华的话又临到我，说：
JER|16|2|“你不可在这地方娶妻，为自己生儿育女。
JER|16|3|因为论到在这地方所生的儿女，又论到在这国中生他们的父母，耶和华如此说：
JER|16|4|他们必死于致命的疾病，无人哀哭，不得埋葬，在地上如粪土，因刀剑和饥荒而灭绝；他们的尸首必给空中的飞鸟和地上的走兽作食物。
JER|16|5|“耶和华如此说：不要进入丧家，不要去哀哭，也不要为他们悲伤，因我已使我的平安、慈爱、怜悯离开这百姓。这是耶和华说的。
JER|16|6|他们连大带小，都必在这地死亡，不得埋葬。人必不为他们哀哭，不为他们割划自己，也不剃光头。
JER|16|7|有丧事，人不为他们擘饼 ，也不因死人安慰他们；他们丧父丧母，人也不给他们一杯酒安慰他们。
JER|16|8|你不可进入宴乐的家，与人同坐又吃又喝，
JER|16|9|因为万军之耶和华－ 以色列 的上帝如此说：看哪，你们还活着的日子，我必在你们眼前止息这地方欢喜和快乐的声音、新郎和新娘的声音。
JER|16|10|“你将这一切的话指示这百姓，他们若问你说：‘耶和华为什么说，要降这大灾祸攻击我们呢？我们有什么罪孽呢？我们向耶和华－我们的上帝犯了什么罪呢？’
JER|16|11|你就对他们说：‘因为你们祖先离弃了我，随从别神，事奉敬拜它们，却离弃我，不遵守我的律法。这是耶和华说的。
JER|16|12|你们行恶比你们祖先更甚，看哪，各人随从自己顽梗的恶心行事，不听从我。
JER|16|13|所以我必将你们从这地赶出，直赶到你们和你们祖先素不认识之地。你们在那里昼夜必事奉别神，因为我必不再向你们施恩。’”
JER|16|14|“看哪，日子将到，人必不再指着那领 以色列 人从 埃及 地上来的永生耶和华起誓。这是耶和华说的。
JER|16|15|人却要指着那领 以色列 人离开北方之地，离开他们被赶到的各国之永生的耶和华起誓；并且我要领他们归回我从前赐给他们祖先之地。”
JER|16|16|“看哪，我要差派许多打鱼的捕获他们；以后，我也要派许多打猎的，从各山上、各冈上、各石穴中猎取他们。这是耶和华说的。
JER|16|17|因我的眼目察看他们一切的行为；他们不能在我面前遮掩，他们的罪孽也不能在我眼前隐藏。
JER|16|18|我要先加倍报应他们的罪孽和罪恶，因为他们以可憎之偶像的尸首使我的地玷污，使我的产业充斥可厌之物。”
JER|16|19|耶和华啊，你是我的力量， 是我的保障， 在患难之日是我的避难所。 列国的人必从地极来到你这里，说： “我们祖先所承受的， 不过是虚假，是虚空无益之物。
JER|16|20|人岂可为自己制造神明呢？ 其实它们不是神明。”
JER|16|21|“所以，看哪，我要使他们知道，就是这一次使他们知道我的手和我的能力。他们就知道我的名是耶和华了。”
JER|17|1|犹大 的罪是用铁笔、用金刚石记录的，铭刻在他们的心版和祭坛角上。
JER|17|2|他们的儿女思念他们在高冈上、青翠树旁的祭坛和 亚舍拉 。
JER|17|3|我田野的山哪，因你在全境内的丘坛所犯的罪，我必使你的财富和一切的财宝成为掠物。
JER|17|4|因自己所做的 ，你必失去我所赐给你的产业。我也必使你在你所不认识的地服侍你的仇敌；因你们激起了我的怒火，直烧到永远。
JER|17|5|耶和华如此说： “倚靠人，以血肉为膀臂， 心中离弃耶和华的， 那人该受诅咒！
JER|17|6|他必像沙漠里的矮树， 不见福乐来到； 他要住在旷野干旱之处， 无人居住的盐地。
JER|17|7|倚靠耶和华、以耶和华为他所仰赖的， 那人有福了！
JER|17|8|他必像树栽于水旁， 在河边扎根， 炎热来到，毫不察觉 ， 叶子仍必青翠； 在干旱之年，一无挂虑， 并且结果不止。
JER|17|9|“人心比万物都诡诈， 坏到极处， 谁能识透呢？
JER|17|10|我－耶和华是鉴察人心，考验人肺腑的， 要按各人所行的和他做事的结果报应他。”
JER|17|11|那不按正道得财富的， 好像鹧鸪孵不是自己生的； 到了中年，财富必离开他， 终久他必成为愚顽人。
JER|17|12|我们的圣所是荣耀的宝座， 从太初就在高处。
JER|17|13|耶和华－ 以色列 的盼望啊， 凡离弃你的必蒙羞。 离我而去的， 他们必被写在地里， 因为他们离弃耶和华，这活水的泉源。
JER|17|14|耶和华啊，求你医治我，我就痊愈， 拯救我，我便得救； 因你是我所赞美的。
JER|17|15|看哪，他们对我说： “耶和华的话在哪里呢？ 让它应验吧！”
JER|17|16|至于我，我并没有逃避作牧人跟随你 ， 也没有想望那灾殃的日子； 这是你所知道的。 我嘴唇所出的都在你面前。
JER|17|17|不要使我因你惊恐； 灾祸来临时，你是我的避难所。
JER|17|18|愿那些迫害我的蒙羞， 却不要使我蒙羞； 使他们惊惶， 却不要使我惊惶； 愿灾祸的日子临到他们， 以加倍的毁坏毁坏他们。
JER|17|19|耶和华对我如此说：“你去站在 犹大 君王出入的 平民门 ，和 耶路撒冷 的各城门口，
JER|17|20|对他们说：‘你们这 犹大 君王、 犹大 众人和 耶路撒冷 所有的居民，凡从这些城门进入的，都当听耶和华的话。
JER|17|21|耶和华如此说：你们要谨慎，不可在安息日挑什么担子进入 耶路撒冷 的城门，
JER|17|22|也不可在安息日从家中挑担子出去。无论何工都不可做，只要以安息日为圣日，正如我所吩咐你们祖先的。’
JER|17|23|他们却不听从，也不侧耳而听，竟硬着颈项不听，不肯领受训诲。
JER|17|24|“你们若留意听从我，在安息日不挑什么担子进入这城的各门，只以安息日为圣日，在那日不做任何工作，这是耶和华说的，
JER|17|25|就必有坐 大卫 宝座的君王和领袖，与 犹大 人，并 耶路撒冷 的居民，或坐车，或骑马，进入这城的各门，而且这城必存到永远。
JER|17|26|也必有人从 犹大 城镇和 耶路撒冷 四围的各处，从 便雅悯 地、 谢非拉 、山区，并 尼革夫 而来，都带燔祭和祭物，素祭和乳香，并感谢祭，到耶和华的殿去。
JER|17|27|你们若不听从我，不以安息日为圣日，仍在安息日挑担子进入 耶路撒冷 的各城门，我必在城门中点火；这火必烧毁 耶路撒冷 的宫殿，不会熄灭。”
JER|18|1|耶和华的话临到 耶利米 ，说：
JER|18|2|“你起来，下到陶匠的家里去，在那里我要使你听见我的话。”
JER|18|3|我就下到陶匠的家里去，看哪，他在转盘上做器皿。
JER|18|4|陶匠用泥做的器皿在他手中做坏了，他就用它另做别的器皿，照他看为好的去做。
JER|18|5|耶和华的话临到我，说：
JER|18|6|“ 以色列 家啊，我待你们岂不能像这陶匠弄泥吗？ 以色列 家，看哪，泥在陶匠的手中怎样，你们在我的手中也怎样。这是耶和华说的。
JER|18|7|我何时论到一邦或一国说，要拔出、拆毁、毁坏；
JER|18|8|我所说的那一邦若回转离开他们的恶，我就改变心意，不将我想要施行的灾祸降与他们。
JER|18|9|我何时论到一邦或一国说，要建立、栽植；
JER|18|10|他们若行我眼中看为恶的事，不听从我的话，我就改变心意，不将我所说的福气赐给他们。
JER|18|11|现在你要对 犹大 人和 耶路撒冷 的居民说：‘耶和华如此说：看哪，我捏塑灾祸降给你们，定意惩罚你们。你们各人当回转离开所行的恶道，改正你们的所作所为。’
JER|18|12|“他们却说：‘没有用的，我们要照自己的计谋去行，各人要随自己顽梗的恶心行事。’”
JER|18|13|“所以，耶和华如此说： 你们且往各国访问， 有谁听见这样的事？ 少女 以色列 行了一件极恐怖的事。
JER|18|14|黎巴嫩 的雪岂能从田野 的磐石上融化呢？ 从远处 流下的凉水岂能干涸呢？
JER|18|15|我的百姓竟忘记我， 向那虚无的神明 烧香， 它们使百姓在所行的路上、在古道上绊跌， 去行未修筑的斜路，
JER|18|16|他们的地就变为荒凉， 长久被人嘲笑； 凡经过这地的必惊骇摇头。
JER|18|17|在仇敌面前，我必如东风刮散他们， 遭难的日子，我要以背向他们， 不以脸看他们。”
JER|18|18|他们说：“来吧！让我们设计谋害 耶利米 ；因为我们有祭司讲律法，有智慧人设谋略，有先知说预言，都未曾断绝。来吧！让我们用舌头攻击他，不要理他一切的话。”
JER|18|19|耶和华啊，求你留心听我， 且听那些指控我的人的话。
JER|18|20|人岂可以恶报善呢？ 他们竟挖坑要害我的性命！ 求你记念我站在你面前为他们说好话， 要使你的愤怒转离他们。
JER|18|21|因此，愿他们的儿女忍受饥荒， 愿他们死于刀剑之手； 愿他们的妻无子，且作寡妇， 愿他们的男人被死亡所灭， 他们的壮丁在阵上被刀击杀。
JER|18|22|你使敌军忽然临到他们的时候， 愿人听见哀声从他们的屋内发出； 因他们挖坑要捉拿我， 暗设罗网要绊我的脚。
JER|18|23|耶和华啊，他们要杀我的那一切计谋， 你都知道。 求你不要赦免他们的罪孽， 也不要从你面前涂去他们的罪恶。 愿他们在你面前跌倒， 愿你在发怒的时候对付他们。
JER|19|1|耶和华如此说：“你去买陶匠的瓷瓶 ，你和 百姓中的长老、位尊的祭司
JER|19|2|出去到 欣嫩子谷 、 哈珥西 的门口，在那里宣告我所吩咐你的话，
JER|19|3|说：‘ 犹大 君王和 耶路撒冷 的居民哪，当听耶和华的话。万军之耶和华－ 以色列 的上帝如此说：看哪，我必使灾祸临到这地方，凡听见的人都必耳鸣；
JER|19|4|因为他们和他们祖先，并 犹大 君王都离弃我，使这地方与我疏远 ，在这里向素不认识的别神烧香，又使这地方遍满无辜人的血。
JER|19|5|他们建造 巴力 的丘坛，要在火中焚烧自己的儿女，作为燔祭献给 巴力 。这不是我命令的，不是我吩咐的，我心里也从来没有想过。
JER|19|6|因此，看哪，日子将到，这地方不再称为 陀斐特 和 欣嫩子谷 ，反倒称为 杀戮谷 。这是耶和华说的。
JER|19|7|我要在这地方使 犹大 和 耶路撒冷 的计谋落空，也必使他们在仇敌面前倒在刀下，倒在寻索其命的人手下。我要把他们的尸首给空中的飞鸟和地上的走兽作食物。
JER|19|8|我必使这城令人惊骇嘲笑；凡路过的，必因这城所遭的灾难惊骇嘲笑。
JER|19|9|仇敌和寻索其命的人追逼他们，使他们落在围困窘迫之中，我必使他们各人吃自己儿女的肉和朋友的肉。’
JER|19|10|“你要在跟你同去的人眼前打碎那瓶，
JER|19|11|对他们说：‘万军之耶和华如此说：我要打碎这百姓和这城，正如人打碎陶匠的器皿，不能再使其完整。他们要在 陀斐特 埋葬，甚至无处可葬。
JER|19|12|我必向这地方和其中的居民如此行，使这城与 陀斐特 一样。这是耶和华说的。
JER|19|13|耶路撒冷 的房屋和 犹大 君王的宫殿，就是他们在其上向天上的万象烧香、向别神献浇酒祭的宫殿房屋，都必被玷污，和 陀斐特 一样。’”
JER|19|14|耶利米 从耶和华差他去说预言的 陀斐特 回来，站在耶和华殿的院中对众百姓说：
JER|19|15|“万军之耶和华－ 以色列 的上帝如此说：‘看哪，我必使我所说的一切灾祸临到这城和属它的城镇，因为他们硬着颈项不听我的话。’”
JER|20|1|音麦 的儿子 巴施户珥 祭司作耶和华殿的总管，听见 耶利米 预言这些事，
JER|20|2|就打 耶利米 先知，用耶和华殿里 上便雅悯门 内的枷锁，把他锁在那里。
JER|20|3|次日， 巴施户珥 开枷释放 耶利米 。于是 耶利米 对他说：“耶和华不叫你的名为 巴施户珥 ，而叫你 玛歌珥．米撒毕 ，
JER|20|4|因耶和华如此说：‘看哪，我要使你和你的众朋友惊吓；你们要亲眼看见他们倒在仇敌的刀下。我必将 犹大 人全都交在 巴比伦 王的手中，他要把他们掳到 巴比伦 去，用刀杀他们。
JER|20|5|我要将这城中一切的货财和劳碌得来的，并一切的珍宝，以及 犹大 君王所有的宝物，都交在仇敌手中。仇敌要抢夺他们，抓住他们，把他们带到 巴比伦 去。
JER|20|6|你， 巴施户珥 ，和所有住在你家中的人都必被掳；你和你的朋友，就是你向他们说假预言的，都要到 巴比伦 去，死在那里，葬在那里。’”
JER|20|7|耶和华啊，你欺哄了我， 我也被你欺哄了。 你比我强，并且得胜。 我终日成为笑柄， 人人都戏弄我。
JER|20|8|我每逢讲话的时候，就哀叹， 我喊叫：“有暴力和毁灭！” 因为耶和华的话终日成了我的凌辱和讥刺。
JER|20|9|我若说：“我不再提耶和华， 也不再奉他的名讲论”， 我心里便觉得 似乎有烧着的火闷在我骨中， 我忍受不住，不能自禁。
JER|20|10|我听见许多的毁谤， 四围都是惊吓； 连我知己朋友都看着我跌倒： “告他吧，我们要告他！ 或者他被引诱， 我们就能胜他， 在他身上报仇。”
JER|20|11|然而，耶和华与我同在， 好像可怕的勇士。 因此，迫害我的都绊跌， 不能得胜； 他们大大蒙羞， 由于行事没有智慧， 必永远受那不能忘怀的羞辱。
JER|20|12|考验义人、察看人肺腑心肠的万军之耶和华啊， 求你使我得见你在他们身上报仇， 因我已将我的案件向你禀明了。
JER|20|13|你们要向耶和华唱歌！ 要赞美耶和华！ 因他救了穷人的性命 脱离恶人的手。
JER|20|14|愿我出生的那日受诅咒！ 愿我母亲生我的那天不蒙福！
JER|20|15|报信给我父亲说 “你得了儿子”， 使我父亲甚欢喜的， 愿那人受诅咒。
JER|20|16|愿那人像耶和华所倾覆而不怜惜的城镇； 愿他早晨听见哀声， 中午听见呐喊；
JER|20|17|因他没有在我未出胎就把我杀了， 以致我母亲成为我的坟墓， 她却一直怀着胎 。
JER|20|18|我为何出胎见劳碌愁苦， 在羞愧中度尽我的年日呢？
JER|21|1|耶和华的话临到 耶利米 。那时， 西底家 王差派 玛基雅 的儿子 巴施户珥 和 玛西雅 的儿子 西番雅 祭司到他那里去，说：
JER|21|2|“请你为我们求问耶和华，因为 巴比伦 王 尼布甲尼撒 前来攻击我们；或者耶和华照他一切奇妙的作为待我们，使 巴比伦 王离开我们而去。”
JER|21|3|耶利米 对他们说：“你们当对 西底家 这样说：
JER|21|4|‘耶和华－ 以色列 的上帝如此说：看哪，我要使你们手中的兵器，就是你们与城外围困你们的 巴比伦 王和 迦勒底 人打仗所用的兵器转回来，把它们聚集在这城中。
JER|21|5|我要在怒气、愤怒和大恼怒中，用伸出来的手和大能的膀臂，亲自攻击你们；
JER|21|6|又要击打这城的居民，他们连人带牲畜都必遭遇大瘟疫而死亡。
JER|21|7|以后，我要将 犹大 王 西底家 和他的臣仆百姓，就是在城内，从瘟疫、刀剑、饥荒中幸存的人，都交在 巴比伦 王 尼布甲尼撒 手中，交在仇敌和寻索其命的人手中。 巴比伦 王必用刀击杀他们，不顾惜，不同情，不怜悯。这是耶和华说的。’
JER|21|8|“你要对这百姓说：‘耶和华如此说：看哪，我将生命的路和死亡的路摆在你们面前。
JER|21|9|住在这城里的必遭刀剑、饥荒、瘟疫而死；但出去投降围困你们之 迦勒底 人的必得存活，保全自己的性命。
JER|21|10|我向这城板脸，降祸不降福；这城必交在 巴比伦 王的手中，他必用火焚烧。这是耶和华说的。’”
JER|21|11|“至于 犹大 王的家，你们当听耶和华的话。
JER|21|12|大卫 家啊，耶和华如此说： ‘每早晨你们要施行公平， 拯救被抢夺的脱离欺压者的手， 免得我的愤怒因你们的恶行发作， 如火燃起，无人能熄灭。’
JER|21|13|住在山谷和平原磐石上的居民啊， 看哪，我与你们为敌， 因为你们说：‘谁能下来攻击我们？ 谁能进入我们的住处呢？’ 这是耶和华说的。
JER|21|14|我必按你们行事的结果惩罚你们， 也必使火在 耶路撒冷 的林中燃起， 将四围所有的尽行烧灭。 这是耶和华说的。”
JER|22|1|耶和华如此说：“你要下到 犹大 王的宫中，在那里说这话，
JER|22|2|你要说：‘坐 大卫 宝座的 犹大 王啊，你和你的臣仆，并进入这些城门的百姓，都当听耶和华的话。
JER|22|3|耶和华如此说：你们要施行公平和公义，拯救被抢夺的脱离欺压者的手，不可亏负寄居的和孤儿寡妇，不可用残暴对待他们，也不可在这地方流无辜人的血。
JER|22|4|你们若切实遵行这话，就必有坐 大卫 宝座的君王和他的臣仆百姓，或坐车或骑马，从这王宫的各门进入。
JER|22|5|你们若不听这些话，我指着自己起誓，这王宫必变为废墟。这是耶和华说的。’
JER|22|6|耶和华论到 犹大 王的家如此说： “我看你如 基列 ， 如 黎巴嫩 的山顶； 然而，我必使你变为旷野， 成为无人居住的城镇。
JER|22|7|我要预备施行毁灭的人， 各人佩带兵器攻击你； 他们要砍伐你佳美的香柏树， 扔在火中。
JER|22|8|“许多国的百姓经过这城，就彼此谈论说：‘耶和华为何向这大城这样做呢？’
JER|22|9|必有人回答说：‘是因他们离弃了耶和华－他们上帝的约，事奉敬拜别神。’”
JER|22|10|不要为已死的人哀哭， 也不要为他悲伤， 却要为离家外出的人大大哀哭； 因为他不再回来见自己的出生地。
JER|22|11|因为论到离开这地方的 约西亚 之子 犹大 王 沙龙 ，就是接续他父亲 约西亚 作王的，耶和华这样说：“他必不再回到这里来，
JER|22|12|却要死在被掳去的地方，必不得再见这地。”
JER|22|13|祸哉！那以不公义盖房，以不公平造楼， 白白使邻舍做工，却不给工钱的人，
JER|22|14|他说：“我要为自己盖宽敞的房，盖高大的楼。” 他为它开窗户， 以香柏木为墙板， 漆上丹红色。
JER|22|15|难道你作王就是要盖香柏木楼房争胜的吗？ 你的父亲岂不是也吃也喝， 也施行公平和公义吗？ 那时他得了福乐。
JER|22|16|他为困苦和贫穷的人伸冤， 那时就得了福乐。 认识我不就在此吗？ 这是耶和华说的。
JER|22|17|你的眼和你的心却专顾不义之财， 流无辜人的血， 行欺压和残暴。
JER|22|18|所以，耶和华论到 约西亚 的儿子 犹大 王 约雅敬 如此说： 人必不为他举哀： “哀哉，我的哥哥！ 哀哉，我的姊姊！” 也不为他举哀： “哀哉，我的主！ 哀哉，我主的荣华！”
JER|22|19|他被埋葬好像埋驴子一样， 被拖出去，扔在 耶路撒冷 城门外。
JER|22|20|你要上 黎巴嫩 哀号， 在 巴珊 扬声， 从 亚巴琳 哀号， 因为你所亲爱的都毁灭了。
JER|22|21|你兴盛的时候，我对你说话； 你却说：“我不听。” 你从年轻时就是这样， 不肯听我的话。
JER|22|22|你的牧人要被风吞吃， 你所亲爱的必被掳去； 那时你必因你一切的恶行抱愧蒙羞。
JER|22|23|你这住 黎巴嫩 、在香柏树上搭窝的， 有痛苦临到你， 如疼痛临到临产的妇人， 那时你何等可怜 ！
JER|22|24|耶和华说：“ 约雅敬 的儿子 犹大 王 哥尼雅 ，虽是我右手上带印的戒指，我凭我的永生起誓，我必将你从其上摘下来。
JER|22|25|我要将你交在寻索你命的人和你所惧怕的人手中，就是 巴比伦 王 尼布甲尼撒 和 迦勒底 人手中。
JER|22|26|我也要将你和生你的母亲赶到别国，不是你们出生的地方；你们必死在那里，
JER|22|27|心中虽然很想归回那地，却不得归回。”
JER|22|28|哥尼雅 这人是被轻看、遭毁坏的罐子， 是无人喜爱的器皿吗？ 他和他的后裔为何被赶到素不认识之地呢？
JER|22|29|地啊，地啊，地啊，当听耶和华的话！
JER|22|30|耶和华如此说： “要把这人登记为无子， 是平生不得亨通的人； 因为他后裔中再无一人得亨通， 能坐在 大卫 的宝座上治理 犹大 。”
JER|23|1|耶和华说：“祸哉！那些残害、赶散我草场之羊的牧人！”
JER|23|2|耶和华－ 以色列 的上帝论到那些牧养他百姓的牧人如此说：“你们赶散我的羊群，并未看顾他们；看哪，我必惩罚你们的恶行。这是耶和华说的。
JER|23|3|我要从我赶他们到的各国召集我羊群中剩余的，领他们归回本处；他们必生养众多。
JER|23|4|我必设立牧人照管他们，牧养他们。他们不再惧怕，不再惊惶，没有一个失丧的。这是耶和华说的。
JER|23|5|“看哪，日子将到，我要为 大卫 兴起公义的苗裔； 他必掌王权，行事有智慧，在地上施行公平和公义。这是耶和华说的。
JER|23|6|在他的日子， 犹大 必得救， 以色列 也安然居住。他的名必称为‘耶和华－我们的义’。
JER|23|7|“看哪，日子将到，人必不再指着那领 以色列 人从 埃及 地上来的永生耶和华起誓。这是耶和华说的。
JER|23|8|人却要指着那领 以色列 家的后裔离开北方之地，离开我赶他们到的各国的永生耶和华起誓。他们必住在本地。”
JER|23|9|论到那些先知， 我心在我里面忧伤， 我的骨头全都发颤； 因耶和华和他的圣言， 我像醉酒的人， 像被酒所胜的人。
JER|23|10|全地满了犯奸淫的人！ 因妄自赌咒，地就悲哀， 旷野的草场都枯干了。 他们所行的道是恶的； 他们的权力用得不对。
JER|23|11|连先知带祭司都是亵渎的， 就是在我殿中，我也看见他们的恶行。 这是耶和华说的。
JER|23|12|因此，他们的道路必像黑暗中的滑地， 他们必被追赶，仆倒在其上； 因为在他们受罚之年， 我必使灾祸临到他们。 这是耶和华说的。
JER|23|13|我在 撒玛利亚 的先知中曾见狂妄的事； 他们藉 巴力 说预言， 使我的百姓 以色列 走迷了路。
JER|23|14|我在 耶路撒冷 的先知中曾见恐怖的事； 他们犯奸淫，行虚谎， 又坚固恶人的手， 无人回转离开自己的恶行。 他们在我面前都像 所多玛 ， 耶路撒冷 的居民都像 蛾摩拉 。
JER|23|15|因此，万军之耶和华论到先知如此说： “看哪，我必使他们吃茵蔯， 喝苦水； 因为亵渎的事出于 耶路撒冷 的先知，遍及各地。”
JER|23|16|万军之耶和华如此说：“你们不要听这些先知向你们所说的预言。他们使你们成为虚无，所说的异象是出于自己的心，不是出于耶和华的口。
JER|23|17|他们常对藐视我的人说：‘耶和华说：你们必享平安。’ 又对一切按自己顽梗之心而行的人说：‘灾祸必不临到你们。’”
JER|23|18|有谁站在耶和华的会中 察看并听见他的话呢？ 有谁留心听他的话呢？
JER|23|19|看哪！耶和华的暴风 在震怒中发出， 是旋转的暴风， 必转到恶人头上。
JER|23|20|耶和华的怒气必不转消， 直到他心中所定的成就了，实现了。 末后的日子，你们要全然明白。
JER|23|21|我并未差遣那些先知， 他们竟自奔跑； 我没有对他们说话， 他们竟自预言。
JER|23|22|他们若站在我的会中， 必使我的百姓听我的话， 又使他们回转离开恶道， 离开他们所行的恶。
JER|23|23|我是靠近你们的上帝，不是遥远的上帝，不是吗？ 这是耶和华说的。
JER|23|24|人岂能在隐密处藏身，使我看不见他呢？这是耶和华说的。我岂不遍满天和地吗？这是耶和华说的。
JER|23|25|我已听见那些先知所说的，他们托我的名说假预言：“我做了梦！我做了梦！”
JER|23|26|所言虚假、心存诡诈的先知，他们这样存心要到几时呢？
JER|23|27|他们彼此述说所做的梦，想要使我的百姓忘记我的名，正如他们祖先因 巴力 忘记我的名一样。
JER|23|28|得梦的先知可以述说那梦；领受我话的人可以诚实讲我的话。糠秕怎能与麦子比较呢？这是耶和华说的。
JER|23|29|我的话岂不像火，又像能打碎磐石的大锤吗？这是耶和华说的。
JER|23|30|看哪，那些先知各从邻舍偷窃我的话，因此我必与他们为敌。这是耶和华说的。
JER|23|31|那些先知用自己的舌头说是耶和华说的；看哪，我必与他们为敌。这是耶和华说的。
JER|23|32|那些以假梦为预言，又述说这梦，以谎言和鲁莽使我百姓走迷了路的，看哪，我必与他们为敌。这是耶和华说的。我并未差遣他们，也没有吩咐他们。他们对这百姓毫无益处。这是耶和华说的。
JER|23|33|无论是这百姓、是先知、是祭司，问你说：“耶和华有什么默示呢？”你就对他们说：“什么默示啊？ 我已撇弃你们了。这是耶和华说的。”
JER|23|34|凡说“耶和华的默示”的，无论是先知、是祭司、是百姓，我必惩罚那人和他的家。
JER|23|35|你们各人要对邻舍、对弟兄如此说：“耶和华回答了什么？耶和华说了什么呢？”
JER|23|36|你们不可再提“耶和华的默示”，因为各人所说的话必成为自己的重担 ；你们错用了永生上帝、万军之耶和华－我们上帝的话。
JER|23|37|你们要对先知如此说：“耶和华回答了你什么？耶和华说了什么呢？”
JER|23|38|你们若说“耶和华的默示”，耶和华就必如此说：“我曾差人到你们那里去，告诉你们不可说‘耶和华的默示’这几个字，你们却说‘耶和华的默示’；
JER|23|39|所以，看哪，我必忘记你们 ，将你们和我所赐给你们并你们祖先的城都撇弃了；
JER|23|40|又必使永远的凌辱和长久的羞耻临到你们，是不能忘记的。”
JER|24|1|巴比伦 王 尼布甲尼撒 将 约雅敬 的儿子 犹大 王 耶哥尼雅 和 犹大 的领袖，并工匠、铁匠从 耶路撒冷 掳去，带到 巴比伦 。这事以后，耶和华指给我看，看哪，有两筐无花果放在耶和华殿前。
JER|24|2|一筐是极好的无花果，像是初熟的；一筐是极坏的无花果，坏得不能吃。
JER|24|3|耶和华对我说：“ 耶利米 ，你看见什么？”我说：“我看见无花果，好的极好，坏的极坏，坏得不能吃。”
JER|24|4|于是耶和华的话临到我，说：
JER|24|5|“耶和华－ 以色列 的上帝如此说：‘被掳去的 犹大 人，就是我所打发离开这地到 迦勒底 人之地去的，我必看顾他们如这好的无花果，使他们得福乐。
JER|24|6|我要眷顾他们，使他们得福乐，领他们归回这地。我也要建立他们，必不拆毁；栽植他们，必不拔出。
JER|24|7|我要赐给他们认识我的心，认识我是耶和华。他们要作我的子民，我要作他们的上帝，他们要一心归向我。’”
JER|24|8|耶和华如此说：“我必将 犹大 王 西底家 和他的众领袖，以及留在这地 耶路撒冷 剩余的人，并住在 埃及 地的 犹大 人都交出来，好像那极坏、坏得不能吃的无花果。
JER|24|9|我必使他们在地上万国中成为恐惧，成为灾祸，在我赶逐他们到的各处成为凌辱、笑柄、讥笑、诅咒的对象。
JER|24|10|我必使刀剑、饥荒、瘟疫临到他们，直到他们从我所赐给他们和他们祖先之地灭绝。”
JER|25|1|约西亚 的儿子 犹大 王 约雅敬 第四年，就是 巴比伦 王 尼布甲尼撒 的元年，耶和华论 犹大 众百姓的话临到 耶利米 。
JER|25|2|耶利米 先知就将这些话对 犹大 众百姓和 耶路撒冷 所有的居民说：
JER|25|3|“从 亚们 的儿子 犹大 王 约西亚 十三年直到今日，在这二十三年中，常有耶和华的话临到我；我也一再对你们传讲，只是你们不听从。
JER|25|4|耶和华也曾一再差遣他的仆人众先知到你们这里来，只是你们不听从，也不侧耳而听，
JER|25|5|说：‘你们各人当回转离开恶道和恶行，就可居住耶和华从古时所赐给你们和你们祖先之地，直到永远。
JER|25|6|不可随从别神，事奉敬拜它们，以你们手所做的惹我发怒；这样，我就不会降灾祸给你们。
JER|25|7|然而你们不听从我，竟以手所做的惹我发怒，害了自己。这是耶和华说的。’”
JER|25|8|所以万军之耶和华如此说：“因为你们不听我的话，
JER|25|9|看哪，我必召北方的众族和我仆人 巴比伦 王 尼布甲尼撒 前来攻击这地和这地的居民，并四围所有的国民。我要将他们尽行灭绝，以致他们令人惊骇、嗤笑，并且永久荒凉 。这是耶和华说的。
JER|25|10|我又要止息他们欢喜和快乐的声音、新郎和新娘的声音、推磨的声音和灯的亮光。
JER|25|11|这全地必然荒凉，令人惊骇。这些国家要服事 巴比伦 王七十年。
JER|25|12|七十年满了以后，我必惩罚 巴比伦 王和那国，并 迦勒底 人之地，因他们的罪孽使那地永远荒凉。这是耶和华说的。
JER|25|13|我也必使我向那地所说的话，就是所有记在这书上， 耶利米 向这些国家说的预言，都临到那地。
JER|25|14|因为必有许多国家和大君王使 迦勒底 人作奴仆；我也必照他们的行为，按他们手所做的报应他们。”
JER|25|15|耶和华－ 以色列 的上帝对我如此说：“你从我手中拿这杯愤怒的酒，给我所差遣你去的各国的百姓喝。
JER|25|16|他们喝了就要东倒西歪，并要发狂，因我使刀剑临到他们中间。”
JER|25|17|我就从耶和华的手中拿了这杯，给耶和华所差遣我去的各国的百姓喝，
JER|25|18|其中有 耶路撒冷 和 犹大 的城镇，并 耶路撒冷 的君王与领袖；因此这城镇荒凉，令人惊骇、嗤笑、诅咒，正如今日一样。
JER|25|19|又有 埃及 王法老和他的臣仆、官长，以及他的众百姓，
JER|25|20|并混居的各族和 乌斯 地的诸王，与 非利士 人之地的诸王，包括 亚实基伦 、 迦萨 、 以革伦 ，以及 亚实突 剩下的人，
JER|25|21|还有 以东 、 摩押 、 亚扪 人，
JER|25|22|推罗 的诸王、 西顿 的诸王、海的那边沿海地区的诸王，
JER|25|23|底但 、 提玛 、 布斯 ，和所有剃鬓发的人，
JER|25|24|阿拉伯 的诸王、住旷野混居各族的诸王、
JER|25|25|心利 的诸王、 以拦 的诸王、 玛代 的诸王、
JER|25|26|北方远近的诸王，以及天下、地面上的万国也一个一个都喝了，以后 示沙克 王也要喝。
JER|25|27|“你要对他们说：‘万军之耶和华－ 以色列 的上帝如此说：你们要喝，且要喝醉，要呕吐，且要跌倒，不再起来，都因我使刀剑临到你们中间。’
JER|25|28|“他们若不肯从你手中拿这杯来喝，你就要对他们说：‘万军之耶和华如此说：你们一定要喝！
JER|25|29|看哪，我既从称为我名下的城起首施行灾祸，你们能免去惩罚吗？你们必不能免，因为我要命刀剑临到地上所有的居民。这是万军之耶和华说的。’
JER|25|30|“所以你要向他们预言这一切的话，对他们说： ‘耶和华从高天吼叫， 从圣所发出声音， 向自己的羊群大声吼叫； 他要向地上所有的居民呐喊， 像踹葡萄的人一样。
JER|25|31|必有响声达到地极， 因为耶和华与列国争辩。 凡有血肉之躯的，他必审问； 至于恶人，他必交给刀剑。 这是耶和华说的。’
JER|25|32|“万军之耶和华如此说： 看哪，必有灾祸发出，从这国到那国， 并有大暴风从地极刮起。
JER|25|33|“到那日，从地这边到地那边，都有耶和华所杀戮的人。必无人哀哭，不得收殓，不得埋葬，必在地面上成为粪土。
JER|25|34|“牧人哪，你们当哀号，呼喊； 羊群的领导者啊，你们要在灰中翻滚； 因为你们被宰杀、被分散 的日子已经来到。 你们要仆倒，好像珍贵的器皿打碎一样。
JER|25|35|牧人无路可逃， 羊群的领导者也无法逃脱。
JER|25|36|听啊，有牧人呼喊， 有羊群领导者哀号的声音， 因为耶和华摧毁他们的草场。
JER|25|37|因耶和华猛烈的怒气， 平安的羊圈都被肃清。
JER|25|38|他像狮子离开洞穴， 他们的地因凶猛的怒气 和他强烈的怒气，都变为荒凉。”
JER|26|1|约西亚 的儿子 犹大 王 约雅敬 登基时，有这话从耶和华临到 耶利米 ，说：
JER|26|2|“耶和华如此说：你要站在耶和华殿的院内，对 犹大 所有城镇的人，就是到耶和华的殿来礼拜的，传讲我所吩咐你的一切话，一字也不可删减。
JER|26|3|或者他们肯听从，各人回转离开恶道，我就改变心意，不将我因他们所行的恶、想要施行的灾祸降与他们。
JER|26|4|你要对他们说，耶和华如此说：‘你们若不听从我，不遵行我在你们面前所设立的律法，
JER|26|5|不听从我一再差遣我仆人众先知到你们那里去所说的话，你们果然没有听从，
JER|26|6|我就必使这殿如 示罗 ，使这城成为地上万国所诅咒的。’”
JER|26|7|耶利米 在耶和华殿中所说的这些话，祭司、先知与众百姓都听见了。
JER|26|8|耶利米 说完了耶和华吩咐他对众百姓说的一切话，祭司、先知与众百姓都来抓住他，说：“你该死！
JER|26|9|你为何假借耶和华的名预言，说这殿必如 示罗 ，这城必荒废无人居住呢？”于是众百姓都聚集在耶和华的殿中围住 耶利米 。
JER|26|10|犹大 的官长们听见这些事，就从王宫上到耶和华的殿，坐在耶和华殿 新门 的入口。
JER|26|11|祭司、先知对官长和众百姓说：“这人该死，因为他说预言攻击这城，正如你们亲耳听见的。”
JER|26|12|耶利米 就对官长和众百姓说：“耶和华差遣我预言攻击这殿和这城，传讲你们所听见的这一切话。
JER|26|13|现在，要改正你们的所作所为，听从耶和华－你们上帝的话，他就必改变心意，不把所说的灾祸降与你们。
JER|26|14|至于我，看哪，我在你们手中，你们眼里看什么是好的，是正确的，就那样待我吧！
JER|26|15|但你们要确实知道，你们若把我处死，就使流无辜人血的罪归给你们和这城，以及城里的居民了；因为耶和华确实差遣我到你们这里来，将这一切话传到你们耳中。”
JER|26|16|官长和众百姓对祭司和先知说：“这人是不该死的，因为他奉耶和华－我们上帝的名向我们说话。”
JER|26|17|国中的长老就有几个人起来，对聚集的众百姓说：
JER|26|18|“当 犹大 王 希西家 的日子，有 摩利沙 人 弥迦 对 犹大 众百姓预言说： ‘万军之耶和华如此说： 锡安 要被耕种像一块田地， 耶路撒冷 要变为废墟， 这殿的山必像丛林的高处。’
JER|26|19|“ 犹大 王 希西家 和 犹大 人岂是把他处死呢？ 希西家 岂不是敬畏耶和华，恳求耶和华施恩吗？耶和华就改变心意，不把所说的灾祸降与他们。若处死这人，我们就做了大恶，害死自己了。”
JER|26|20|有一个人，就是 示玛雅 的儿子 基列．耶琳 人 乌利亚 ，也奉耶和华的名说预言；他说预言攻击这城和这地，和 耶利米 所说的完全一样。
JER|26|21|约雅敬 王和他所有的勇士、官长听见了 乌利亚 的话，王想要把他处死。 乌利亚 听见就惧怕，逃往 埃及 去了。
JER|26|22|约雅敬 王差 亚革波 的儿子 以利拿单 ，带领几个人前往 埃及 。
JER|26|23|他们将 乌利亚 从 埃及 带出来，解送到 约雅敬 王那里；王用刀杀了他，把他的尸首抛在平民的坟地中。
JER|26|24|然而， 沙番 的儿子 亚希甘 保护 耶利米 ，不将他交在百姓手中，以免他们把他处死。
JER|27|1|约西亚 的儿子 犹大 王 约雅敬 登基时，有这话从耶和华临到 耶利米 ，说：
JER|27|2|“耶和华对我如此说：你要为自己做皮带和木轭，套在你的颈项上，
JER|27|3|然后托那些来到 耶路撒冷 ，到 犹大 王 西底家 那里的使节，把皮带和木轭送到 以东 王、 摩押 王、 亚扪 王、 推罗 王、 西顿 王那里，
JER|27|4|且嘱咐他们转达他们的主人。万军之耶和华－ 以色列 的上帝如此说，你们要对你们的主人这样说：
JER|27|5|我用大能和伸出来的膀臂创造大地和地上的人民、牲畜。我看给谁合适，就把地给谁。
JER|27|6|现在我将全地都交在我仆人 巴比伦 王 尼布甲尼撒 手中，也把野地的走兽给他使用。
JER|27|7|列国都要服事他和他的子孙，直到他本国遭报的日期来到；那时，许多国家和大君王要使他作奴隶。
JER|27|8|“无论哪一邦、哪一国，不肯服事 巴比伦 王 尼布甲尼撒 ，不把颈项放在他的轭下，我必用刀剑、饥荒、瘟疫惩罚那邦，直到我藉 巴比伦 王的手毁灭他们。这是耶和华说的。
JER|27|9|至于你们，不可听从你们的先知和占卜的、做梦的 、观星象的，以及行邪术的；他们对你们说：‘你们必不致服事 巴比伦 王。’
JER|27|10|他们向你们传的是假预言，要叫你们远离本地，以致我将你们赶出去，使你们灭亡。
JER|27|11|但哪一邦肯把颈项放在 巴比伦 王的轭下服事他，我必使那邦仍在本地存留，在那里耕种居住。这是耶和华说的。”
JER|27|12|我就照这一切话对犹大王 西底家 说：“你们要把颈项放在 巴比伦 王的轭下，服事他和他的百姓，就得存活。
JER|27|13|你和你的百姓何必因刀剑、饥荒、瘟疫而死亡，像耶和华所论不肯服事 巴比伦 王的国家呢？
JER|27|14|不可听那些先知对你们所说的话，他们说：‘你们必不致服事 巴比伦 王’，其实他们向你们传的是假预言。
JER|27|15|耶和华说：‘我并未差遣他们，他们却托我的名传假预言，使我将你们和向你们说预言的那些先知赶出去，一同灭亡。’”
JER|27|16|我又对祭司和这众百姓说：“耶和华如此说：你们不可听那先知对你们所说的预言，他们说：‘看哪，耶和华殿中的器皿快要从 巴比伦 带回来’；其实他们向你们传的是假预言。
JER|27|17|不可听从他们，只管服事 巴比伦 王，就得存活。何必使这城变为废墟呢？
JER|27|18|他们若真是先知，有耶和华的话临到他们，让他们祈求万军之耶和华，使耶和华殿中和 犹大 王宫内，并 耶路撒冷 剩下的器皿，不致被带到 巴比伦 去。
JER|27|19|万军之耶和华这样论柱子、铜海、盆座，并留在这城里剩下的器皿，
JER|27|20|就是 巴比伦 王 尼布甲尼撒 掳掠 约雅敬 的儿子 犹大 王 耶哥尼雅 ，并 犹大 、 耶路撒冷 所有贵族时，没有从 耶路撒冷 掠去 巴比伦 的器皿。
JER|27|21|论到那在耶和华殿中和 犹大 王宫内，并 耶路撒冷 剩下的器皿，万军之耶和华－ 以色列 的上帝如此说：
JER|27|22|它们必被带到 巴比伦 ，存放在那里，直到我眷顾 以色列 人，将这些器皿带回归还此地的日子。这是耶和华说的。”
JER|28|1|当年，就是 犹大 王 西底家 登基第四年五月， 押朔 的儿子 基遍 人 哈拿尼雅 先知，在耶和华的殿中当着祭司和众百姓的面对我说：
JER|28|2|“万军之耶和华－ 以色列 的上帝如此说：我已经折断 巴比伦 王的轭。
JER|28|3|二年之内，我要将 巴比伦 王 尼布甲尼撒 从这地掳掠到 巴比伦 的器皿，就是耶和华殿中的一切器皿，都带回此地。
JER|28|4|我又要将 约雅敬 的儿子 犹大 王 耶哥尼雅 和被掳到 巴比伦 所有的 犹大 人带回此地，因为我要折断 巴比伦 王的轭。这是耶和华说的。”
JER|28|5|耶利米 先知当着祭司和站在耶和华殿里众百姓的面，对 哈拿尼雅 先知说：
JER|28|6|“阿们！愿耶和华如此行，愿耶和华实现你所预言的话，将耶和华殿中的器皿和所有被掳去的人从 巴比伦 带回此地。
JER|28|7|然而我在你和众百姓耳中所要说的话，你应当听。
JER|28|8|从古以来，在你我以前的众先知，向多国和大邦说预言，论到战争、灾祸 、瘟疫的事。
JER|28|9|至于那预言平安的先知，到先知的话应验的时候，人就知道他真是耶和华所差来的。”
JER|28|10|哈拿尼雅 先知就取下 耶利米 先知颈项上的轭，把它折断。
JER|28|11|哈拿尼雅 又当着众百姓的面说：“耶和华如此说：二年之内我必照样从列国的颈项上折断 巴比伦 王 尼布甲尼撒 的轭。” 耶利米 先知就离开了。
JER|28|12|哈拿尼雅 先知折断 耶利米 先知颈项上的轭以后，耶和华的话临到 耶利米 ，说：
JER|28|13|“你去告诉 哈拿尼雅 说，耶和华如此说：你折断木轭，却换来铁轭！
JER|28|14|万军之耶和华－ 以色列 的上帝如此说：我已将铁轭加在这些国的颈项上，使他们服事 巴比伦 王 尼布甲尼撒 。他们总要服事他，我也把野地的走兽给了他。”
JER|28|15|于是 耶利米 先知对 哈拿尼雅 先知说：“ 哈拿尼雅 啊，你应当听！耶和华并没有差遣你，你竟使这百姓倚靠谎言。
JER|28|16|所以耶和华如此说：看哪，我要把你从地面上除掉，你今年必死，因为你向耶和华说了叛逆的话。”
JER|28|17|这样， 哈拿尼雅 先知当年七月间就死了。
JER|29|1|耶利米 先知从 耶路撒冷 送信给被掳幸存的长老，以及祭司、先知，和 尼布甲尼撒 从 耶路撒冷 掳到 巴比伦 去的众百姓。
JER|29|2|这是在 耶哥尼雅 王和太后、官员，并 犹大 和 耶路撒冷 的领袖，以及工匠、铁匠都离开 耶路撒冷 之后。
JER|29|3|他藉 沙番 的儿子 以利亚萨 和 希勒家 的儿子 基玛利 的手送去；他们二人是 犹大 王 西底家 差往 巴比伦 去见 巴比伦 王 尼布甲尼撒 的。
JER|29|4|信上说：“万军之耶和华－ 以色列 的上帝对所有被掳的，就是我使他们从 耶路撒冷 被掳到 巴比伦 去的人如此说：
JER|29|5|你们要建造房屋，住在其中；要开垦田园，吃园中所出产的；
JER|29|6|要娶妻生儿养女，为你们的儿子娶妻，使你们的女儿嫁人，生儿养女。你们要在那里生养众多，不可减少。
JER|29|7|我使你们被掳到的那城，你们要为那城求平安，为那城向耶和华祈求，因为那城得平安，你们也随着得平安。
JER|29|8|万军之耶和华－ 以色列 的上帝如此说：不要被你们中间的先知和占卜的所诱惑，也不要听信你们 所做的梦，
JER|29|9|因为他们托我的名对你们说假预言，我并未差遣他们。这是耶和华说的。
JER|29|10|“耶和华如此说：为 巴比伦 所定的七十年满了以后，我要眷顾你们，向你们实现我的恩言，使你们归回此地。
JER|29|11|我知道我向你们所怀的意念是赐平安的意念，不是降灾祸的意念，要叫你们末后有指望。这是耶和华说的。
JER|29|12|你们呼求我，向我祷告，我就应允你们。
JER|29|13|你们寻求我，若专心寻求我，就必寻见。
JER|29|14|我必被你们寻见，也必使你们被掳的人归回。这是耶和华说的。我必将你们从各国和我赶你们到的各处召集过来，又将你们带回我使你们被掳离开的地方。这是耶和华说的。
JER|29|15|“你们说：‘耶和华已在 巴比伦 为我们兴起先知。’
JER|29|16|所以耶和华如此论坐 大卫 宝座的君王和住在这城里所有的百姓，就是未曾与你们一同被掳的弟兄，
JER|29|17|万军之耶和华如此说：‘看哪，我必使刀剑、饥荒、瘟疫临到他们，使他们像极坏的无花果，坏得不能吃。
JER|29|18|我必用刀剑、饥荒、瘟疫追赶他们，使地上万国因他们而惊骇；在我赶他们到的各国，令人诅咒、惊骇、嗤笑、羞辱。
JER|29|19|这是因为他们不听从我先前一再差遣我仆人众先知说的话。这是耶和华说的。你们 也一样不听。这是耶和华说的。’
JER|29|20|所以你们所有被掳去的，就是我从 耶路撒冷 放逐到 巴比伦 去的，当听耶和华的话。
JER|29|21|万军之耶和华－ 以色列 的上帝论 哥赖雅 的儿子 亚哈 和 玛西雅 的儿子 西底家 如此说：‘他们托我的名向你们说假预言，看哪，我必把他们交在 巴比伦 王 尼布甲尼撒 的手中，他要在你们眼前杀害他们。
JER|29|22|在 巴比伦 所有被掳的 犹大 人必藉这二人赌咒说：愿耶和华使你像 巴比伦 王在火中焚烧的 西底家 和 亚哈 一样。
JER|29|23|这二人在 以色列 中做了丑事，与邻舍的妻行淫，又假托我的名说我未曾吩咐他们的话。我知道这一切，也作见证。这是耶和华说的。’”
JER|29|24|“你要对 尼希兰 人 示玛雅 说：
JER|29|25|万军之耶和华－ 以色列 的上帝如此说：你曾用自己的名送信给 耶路撒冷 的众百姓和 玛西雅 的儿子 西番雅 祭司，并众祭司，说：
JER|29|26|‘耶和华已经立你 西番雅 为祭司，代替 耶何耶大 祭司，使耶和华的殿中有总管，好把所有狂妄自称先知的人用枷枷住，用锁锁住。
JER|29|27|现在 亚拿突 人 耶利米 向你们自称先知，你为什么不责备他呢？
JER|29|28|他送信给我们在 巴比伦 的人说：被掳的事必长久，你们要建造房屋，住在其中；要开垦田园，吃园中所出产的。’”
JER|29|29|西番雅 祭司就把这信念给 耶利米 先知听。
JER|29|30|于是耶和华的话临到 耶利米 ，说：
JER|29|31|“你当送信给所有被掳的人，说：‘耶和华论到 尼希兰 人 示玛雅 说：因为 示玛雅 向你们说预言，使你们倚靠谎言，而我并没有差遣他，
JER|29|32|所以耶和华如此说：看哪，我必惩罚 尼希兰 人 示玛雅 和他的后裔，他必无一人存留住在这民中，也看不见我所要赏赐给我百姓的福乐，因为他向耶和华说了叛逆的话。这是耶和华说的。’”
JER|30|1|耶和华的话临到 耶利米 ，说：
JER|30|2|“耶和华－ 以色列 的上帝如此说：你要将我对你说过的一切话都写在书上。
JER|30|3|看哪，日子将到，我要使我的百姓 以色列 和 犹大 被掳的人归回。这是耶和华说的。耶和华说：我要使他们回到我所赐给他们祖先之地，他们就得这地为业。”
JER|30|4|以下是耶和华论到 以色列 和 犹大 所说的话：
JER|30|5|耶和华如此说： “我们听见颤抖的声音， 令人惧怕，没有平安。
JER|30|6|你们且访查看看， 男人会生孩子吗？ 我怎么看见人人都用手撑腰， 像临产的妇人， 脸都发白了呢？
JER|30|7|哀哉！ 那日为大， 无日可比； 这是 雅各 遭难的时刻， 但他必从患难中得拯救。”
JER|30|8|万军之耶和华说：“到那日，我必折断你颈项上仇敌的轭，拉断你的皮带。陌生人必不再使他作奴隶。
JER|30|9|他们却要事奉耶和华－他们的上帝，事奉我为他们所兴起的 大卫 王。”
JER|30|10|我的仆人 雅各 啊，不要惧怕； 以色列 啊，不要惊惶； 因我从远方拯救你， 从被掳之地拯救你的后裔； 雅各 必回来得享平静安逸， 无人能使他害怕。 这是耶和华说的。
JER|30|11|因我与你同在，要拯救你， 也要将那些国灭绝净尽， 就是我赶你去的那些国； 却不将你灭绝净尽， 倒要从宽惩治你， 但绝不能不罚你。 这是耶和华说的。
JER|30|12|耶和华如此说： “你的损伤无法医治， 你的伤痕极其重大。
JER|30|13|无人为你的伤痛辩护， 也没有可医治你的良药。
JER|30|14|你所亲爱的都忘记你， 不来探望你。 我因你罪孽甚大，罪恶众多， 曾藉仇敌加的伤害伤害你， 藉残忍者惩治你。
JER|30|15|你为何因所受的损伤哀号呢？ 你的痛苦无法医治。 我因你罪孽甚大，罪恶众多， 曾将这些加在你身上。
JER|30|16|因此，凡吞吃你的必被吞吃， 你的敌人个个都被掳去； 掳掠你的必成为掳物， 我使抢夺你的成为掠物。
JER|30|17|我必使你痊愈， 医好你的伤痕， 都因人称你为被赶散的， 这是 锡安 ，是无人来探望的！ 这是耶和华说的。”
JER|30|18|耶和华如此说： “看哪，我必使 雅各 被掳去的帐棚归回， 也必顾惜他的住处。 城必建造在原有的废墟上， 宫殿也必照样有人居住。
JER|30|19|必有感谢和欢乐的声音从其中发出， 我使他们增多，不致减少； 使他们尊荣，不致卑微。
JER|30|20|他们的儿女必如往昔； 他们的会众坚立在我面前； 凡欺压他们的，我必惩罚。
JER|30|21|他们的君王是他们自己的人， 掌权的必出自他们。 我要使他接近我， 他也要亲近我； 不然，谁敢放胆亲近我呢？ 这是耶和华说的。
JER|30|22|你们要作我的子民， 我要作你们的上帝。”
JER|30|23|看哪，耶和华的愤怒 如暴风已经发出； 是扫灭的暴风， 必转到恶人的头上。
JER|30|24|耶和华的烈怒必不转消， 直到他心中所定的成就了，实现了； 末后的日子你们就会明白。
JER|31|1|耶和华说：“那时，我必作 以色列 各家的上帝，他们必作我的子民。”
JER|31|2|耶和华如此说： “从刀剑生还的百姓 在旷野蒙恩； 以色列 寻找安歇之处。”
JER|31|3|耶和华从远方向我显现： “我以永远的爱爱你， 因此，我以慈爱吸引你。”
JER|31|4|少女 以色列 啊， 我要再建立你，你就得以建立； 你必再拿起手鼓， 随着欢乐的舞者而出。
JER|31|5|你必在 撒玛利亚 的山上栽葡萄园， 栽种的人栽种，而且享用。
JER|31|6|日子将到，守望的人必在 以法莲 山上呼叫： “起来吧！我们要上 锡安 ， 到耶和华－我们的上帝那里去。”
JER|31|7|耶和华如此说： “你们当为 雅各 欢乐歌唱， 为万国中为首的欢呼。 当传扬，颂赞说： ‘耶和华啊， 求你拯救你的百姓 ， 拯救 以色列 的余民。’
JER|31|8|看哪，我必将他们从北方之地领来， 从地极召集而来； 同他们来的有盲人、瘸子、孕妇、产妇； 他们必成群结队回到这里。
JER|31|9|他们要哭泣而来。 我要照他们恳求的引导他们， 使他们在河水旁行走正直的路， 他们在其上必不致绊跌； 因为我是 以色列 的父， 以法莲 是我的长子。
JER|31|10|列国啊，要听耶和华的话， 要在远方的海岛传扬，说： “赶散 以色列 的必召集他， 看守他，如牧人看守羊群。”
JER|31|11|因为耶和华救赎了 雅各 ， 救赎他脱离比他更强之人的手。
JER|31|12|他们来到 锡安 的高处歌唱， 因耶和华的宏恩而喜乐洋溢， 就是五谷、新酒和新的油， 并羔羊和牛犊。 他们必像有水浇灌的园子， 一点也不再有愁烦。
JER|31|13|那时，少女必欢乐跳舞； 年轻的、年老的，都一同欢乐； 因为我要使他们的悲哀变为欢喜， 并要安慰他们，使他们的愁烦转为喜乐。
JER|31|14|我必以肥油使祭司的心满足， 我的百姓也要因我的恩惠知足。 这是耶和华说的。
JER|31|15|耶和华如此说： “在 拉玛 听见号啕痛哭的声音， 是 拉结 哭她儿女，不肯因她儿女受安慰， 因为他们都不在了。”
JER|31|16|耶和华如此说： “不要出声哀哭， 你的眼目也不要流泪； 因你的辛劳必有报偿， 他们必从仇敌之地归回。 这是耶和华说的。
JER|31|17|你末后必有指望， 你的儿女必回到自己的疆土。 这是耶和华说的。
JER|31|18|我听见 以法莲 为自己悲叹说： ‘你管教我，我便受管教， 我如未驯服的牛犊。 求你使我回转，我便回转， 因为你是耶和华－我的上帝。
JER|31|19|我背离以后就懊悔， 受教以后就捶胸 ； 我因担当年轻时的凌辱就抱愧蒙羞。’
JER|31|20|以法莲 是我的爱子吗？ 是我喜欢的孩子吗？ 我每逢责备他，仍深顾念他。 因此，我的心肠牵挂着他， 我必要怜悯他。 这是耶和华说的。
JER|31|21|少女 以色列 啊， 当为自己设立路标， 为自己竖起指路牌。 要留心向着大道， 就是你曾走过的路； 你当回转，回到你自己的城镇。
JER|31|22|背道的女子啊， 你翻来覆去要到几时呢？ 耶和华在地上造了一件新事， 就是女子护卫男子。”
JER|31|23|万军之耶和华－ 以色列 的上帝如此说：“我使被掳之人归回的时候，他们在 犹大 地和其中的城镇必再这样说： 公义的居所啊，圣山哪， 愿耶和华赐福给你。
JER|31|24|犹大 和 犹大 城镇的人，耕地的和带着群畜游牧的人，都要一同住在其中。
JER|31|25|疲乏的人，我使他振作；愁烦的人，我使他满足。”
JER|31|26|于是我醒了，我看到我睡得香甜。
JER|31|27|“看哪，日子将到，我要使人的后代和牲畜的种，在 以色列 家和 犹大 家繁衍。这是耶和华说的。
JER|31|28|我先前怎样看守他们，为要拔出、拆毁、毁坏、倾覆、苦害，也必照样看守他们，为要建立、栽植。这是耶和华说的。
JER|31|29|当那些日子，人不再说： ‘父亲吃了酸葡萄， 儿子牙齿就酸倒。’
JER|31|30|但各人要因自己的罪死亡；凡吃酸葡萄的，自己的牙必酸倒。
JER|31|31|“看哪，日子将到，我要与 以色列 家和 犹大 家另立新的约。这是耶和华说的。
JER|31|32|这约不像我拉着他们祖宗的手，领他们出 埃及 地的时候与他们所立的约。我虽作他们的丈夫，他们却背了我的约。这是耶和华说的。
JER|31|33|那些日子以后，我与 以色列 家所立的约是这样：我要将我的律法放在他们里面，写在他们心上。我要作他们的上帝，他们要作我的子民。这是耶和华说的。
JER|31|34|他们各人不再教导自己的邻舍和弟兄说：‘你该认识耶和华’，因为他们从最小的到最大的都必认识我。我要赦免他们的罪孽，不再记得他们的罪恶。这是耶和华说的。”
JER|31|35|耶和华使太阳白昼发光， 按定例使月亮和星辰照耀黑夜， 又搅动大海，使海中波浪澎湃， 万军之耶和华是他的名， 他如此说：
JER|31|36|“这些定例若能在我面前废掉， 以色列 的后裔才会在我面前断绝， 永远不再成国。 这是耶和华说的。”
JER|31|37|耶和华如此说： “若有人能测量上面的天， 探索下面地的根基， 我才会因 以色列 后裔所做的一切弃绝他们。 这是耶和华说的。”
JER|31|38|看哪，日子将到，这城必为耶和华而造，从 哈楠业楼 直到 角门 。这是耶和华说的。
JER|31|39|丈量的绳子要往外拉出，直到 迦立山 ，又转到 歌亚 ；
JER|31|40|抛尸的全谷和倒灰之处，并一切田地，直到 汲沦溪 ，又到东边 马门 的角落，都要归耶和华为圣；不再拔出，不再倾覆，直到永远。
JER|32|1|犹大 王 西底家 第十年，就是 尼布甲尼撒 十八年，耶和华的话临到 耶利米 。
JER|32|2|那时 巴比伦 王的军队围困 耶路撒冷 ， 耶利米 先知被囚在 犹大 王宫中护卫兵的院内；
JER|32|3|因为 犹大 王 西底家 囚禁他，说：“你为什么预言耶和华如此说：‘看哪，我要把这城交在 巴比伦 王的手中，他必攻下这城。
JER|32|4|犹大 王 西底家 必不能逃脱 迦勒底 人的手，定要交在 巴比伦 王手中，他要亲眼看到 巴比伦 王，亲口跟他说话。
JER|32|5|巴比伦 王要将 西底家 带到 巴比伦 ； 西底家 必住在那里，直到我惩罚 他的时候。你们虽与 迦勒底 人争战，却不顺利。这是耶和华说的。’”
JER|32|6|耶利米 说：“耶和华的话临到我，说：
JER|32|7|‘看哪，你叔父 沙龙 的儿子 哈拿篾 必到你这里来，说：请你买我在 亚拿突 的那块地，因为你有代赎的责任。’
JER|32|8|我叔父的儿子 哈拿篾 果然照耶和华的话来到护卫兵的院内，对我说：‘请你买我在 便雅悯 境内、 亚拿突 的那块地；因为它应该由你来承受，而且你也有代赎的责任。请你买下它吧！’我就知道这确是耶和华的话。
JER|32|9|“我便向我叔父的儿子 哈拿篾 买了 亚拿突 的那块地，秤了十七舍客勒银子给他。
JER|32|10|我在契上签字，将契封缄，又请证人来，用天平把银子秤给他。
JER|32|11|我又将按照法定条例所立的买契，就是封缄的那一张和敞开的那一张，
JER|32|12|在我叔父的儿子 哈拿篾 和签字作证的人，并坐在护卫兵院内所有 犹大 人眼前，交给 玛西雅 的孙子 尼利亚 的儿子 巴录 。
JER|32|13|我在众人眼前嘱咐 巴录 说：
JER|32|14|‘万军之耶和华－ 以色列 的上帝如此说：你拿着这文件，就是封缄的和敞开的买契，把它们放在瓦器里，以便长久保存。
JER|32|15|因为万军之耶和华－ 以色列 的上帝如此说：将来在这地必有人再购置房屋、田地和葡萄园。’”
JER|32|16|“我将买契交给 尼利亚 的儿子 巴录 以后，就向耶和华祷告说：
JER|32|17|‘唉！主耶和华，看哪，你曾用大能和伸出来的膀臂创造天和地，在你没有难成的事。
JER|32|18|你施慈爱给千万人，又将祖先的罪孽报应在他后世子孙身上。至大全能的上帝啊，万军之耶和华是你的名，
JER|32|19|你谋事有大略，行事有大能，注目观看世人一切的举动，为要照各人所做的和他做事的结果报应他。
JER|32|20|你在 埃及 地显神迹奇事，直到今日在 以色列 和世人中间也是如此，建立了自己的名声，正如今日一样。
JER|32|21|你用神迹奇事、大能的手、伸出来的膀臂和大可畏的事，领你的百姓 以色列 出了 埃及 ，
JER|32|22|把这地赏赐给他们，就是你向他们列祖起誓应许要赐给他们的流奶与蜜之地。
JER|32|23|他们进入并取得这地，却不听从你的话，也不遵行你的律法。你吩咐他们所当行的，他们都不去行，因此你使这一切的灾祸临到他们。
JER|32|24|看哪，敌人已经来到，用土堆攻取这城；这城也因刀剑、饥荒、瘟疫被交在攻城的 迦勒底 人手中。你所说的话都应验了，看哪，你也看见了。
JER|32|25|主耶和华啊，你却对我说，要用银子为自己买那块地，又请人作证；其实这城已交在 迦勒底 人的手中了。’”
JER|32|26|耶和华的话临到 耶利米 ，说：
JER|32|27|“看哪，我是耶和华，是凡有血肉之躯者的上帝，在我岂有难成的事吗？
JER|32|28|耶和华如此说：看哪，我必将这城交给 迦勒底 人的手和 巴比伦 王 尼布甲尼撒 的手，他必攻取这城。
JER|32|29|攻城的 迦勒底 人必来放火焚烧这城和城里的房屋；人曾在这房顶上向 巴力 烧香，向别神献浇酒祭，惹我发怒。
JER|32|30|以色列 人和 犹大 人从年轻时，就专做我眼中看为恶的事。 以色列 人尽以手所做的惹我发怒。这是耶和华说的。
JER|32|31|这城自从建造的那日直到今日，常惹我的怒气和愤怒，以致我将这城从我面前除掉；
JER|32|32|这是因 以色列 人和 犹大 人一切的邪恶，就是他们和他们的君王、官长、祭司、先知，并 犹大 人，以及 耶路撒冷 居民所做的，惹我发怒。
JER|32|33|他们以背向我，不以面向我；我虽然一再教导他们，他们却不听从，不领受训诲，
JER|32|34|竟把可憎之偶像设立在称为我名下的殿中，玷污了这殿。
JER|32|35|他们在 欣嫩子谷 建造 巴力 的丘坛，把自己的儿女经火献给 摩洛 ；他们行这可憎的事，使 犹大 陷在罪里，这并不是我吩咐的，我心里也从来没有想过。”
JER|32|36|现在论到这城，就是你们所说，已经因刀剑、饥荒、瘟疫被交在 巴比伦 王手中的，耶和华－ 以色列 的上帝如此说：
JER|32|37|“看哪，我曾在怒气、愤怒和大恼怒中，将 以色列 人赶到各国；我必从那里将他们召集出来，领他们回到此地，使他们安然居住。
JER|32|38|他们要作我的子民，我要作他们的上帝。
JER|32|39|我要使他们彼此同心同道，好叫他们永远敬畏我，使他们和他们后世的子孙得享福乐。
JER|32|40|我要跟他们立永远的约，要施恩给他们，绝不转离；又要把敬畏我的心放在他们心里，不离弃我。
JER|32|41|我必欢喜施恩给他们，尽心尽意、真诚地将他们栽于此地。
JER|32|42|“因为耶和华如此说：我怎样使这一切大灾祸临到这百姓，也要照样使我所应许他们的一切福乐都临到他们。
JER|32|43|你们所说荒凉、无人、无牲畜，已交给 迦勒底 人手的这地，必有人购置田地。
JER|32|44|在 便雅悯 地、 耶路撒冷 四围的各处、 犹大 的城镇、山区的城镇、 谢非拉 的城镇，并 尼革夫 的城镇，人必用银子买田地，在契上签字，将契封缄，找人作证，因为我必使被掳的人归回。这是耶和华说的。”
JER|33|1|耶利米 还囚在护卫兵的院内，耶和华的话第二次临到他，说：
JER|33|2|“成事的耶和华，塑造它为要建立它的耶和华，名为耶和华的那位如此说：
JER|33|3|‘你求告我，我就应允你，并将你所不知道、又大又隐密的事指示你。
JER|33|4|论到这城中的房屋和 犹大 君王的宫殿，就是拆毁来挡围城工事和刀剑的，耶和华－ 以色列 的上帝如此说：
JER|33|5|他们与 迦勒底 人争战，用我在怒气和愤怒中所杀之人的尸首塞满这房屋；我因他们一切的恶，转脸不顾这城。
JER|33|6|看哪，我要使这城得以痊愈安舒，我要医治他们，将丰盛的平安与信实显明给他们。
JER|33|7|我也要使 犹大 被掳的和 以色列 被掳的人归回，并要建立他们，如起初一样。
JER|33|8|我要洗净他们干犯我的一切罪，赦免他们干犯我、违背我的一切罪。
JER|33|9|这城在地上万国面前要因我的缘故，以喜乐得名，得颂赞，得荣耀，因为他们听见我所赏赐的一切福乐。他们因我向这城所施的一切福乐平安，就惧怕战兢。”
JER|33|10|耶和华如此说：“你们论这地方，说是荒废、无人、无牲畜之地，但在这荒凉、无人、无居民、无牲畜的 犹大 城镇和 耶路撒冷 街上，必再听见
JER|33|11|欢喜和快乐的声音、新郎和新娘的声音，并听见有人说： 你们要称谢万军之耶和华， 因耶和华本为善， 他的慈爱永远长存！ 他们奉感谢祭到耶和华的殿中；因为我必使这地被掳的人归回，如起初一样。这是耶和华说的。”
JER|33|12|万军之耶和华如此说：“在这荒废、无人、无牲畜之地，并其中所有的城镇，必再有牧人的草场，可让羊群躺卧在那里。
JER|33|13|在山区的城镇、 谢非拉 的城镇、 尼革夫 的城镇、 便雅悯 地、 耶路撒冷 四围的各处和 犹大 的城镇，必再有羊群从数点的人手下经过。这是耶和华说的。
JER|33|14|“看哪，日子将到，我应许 以色列 家和 犹大 家的恩言必然实现。这是耶和华说的。
JER|33|15|在那些日子、那时候，我必使 大卫 公义的苗裔长起来；他必在地上施行公平和公义。
JER|33|16|在那些日子， 犹大 必得救， 耶路撒冷 必安然居住，他的名必称为‘耶和华－我们的义’。
JER|33|17|“因为耶和华如此说： 大卫 家必永远不断有人坐在 以色列 家的宝座上；
JER|33|18|利未 家的祭司也不断有人在我面前献燔祭、烧素祭，时常办理献祭的事。”
JER|33|19|耶和华的话临到 耶利米 ，说：
JER|33|20|“耶和华如此说：你们若能废弃我所立白日黑夜的约，使白日黑夜不按时轮转，
JER|33|21|就能废弃我与我仆人 大卫 所立的约，使他没有后裔在他的宝座上作王，并能废弃我与事奉我的 利未 家的祭司所立的约。
JER|33|22|正如天上的万象不能数算，海边的尘沙不能斗量，我必照样使我仆人 大卫 的后裔和事奉我的 利未 人多起来。”
JER|33|23|耶和华的话临到 耶利米 ，说：
JER|33|24|“你没有留意这百姓所说的话吗？他们说：‘耶和华所拣选的二族，他已经弃绝了。’他们这样藐视我的百姓，不把他们当作国来看待。
JER|33|25|耶和华如此说：除非我没有立白日黑夜之约，也未曾安排天和地的定例，
JER|33|26|否则我不会弃绝 雅各 的后裔和我仆人 大卫 的后裔，使 大卫 的后裔不再治理 亚伯拉罕 、 以撒 、 雅各 的后裔。我必使他们被掳的人归回，也必怜悯他们。”
JER|34|1|巴比伦 王 尼布甲尼撒 率领他的全军和地上他管辖的各国各邦，攻打 耶路撒冷 和 耶路撒冷 所有的城镇。那时，耶和华的话临到 耶利米 ，说：
JER|34|2|“耶和华－ 以色列 的上帝说，你去告诉 犹大 王 西底家 ，耶和华如此说：看哪，我要把这城交在 巴比伦 王的手中，他必用火焚烧。
JER|34|3|你必不能逃脱他的手，定被拿住，交在他手中。你要亲眼看到 巴比伦 王，他要亲口跟你说话，你也必到 巴比伦 去。
JER|34|4|犹大 王 西底家 啊，你一定要听耶和华的话。耶和华论到你如此说：你必不死于刀下；
JER|34|5|必平安而终，人要为你焚烧，好像为你祖先，就是在你以前早先的王焚烧一样。人要为你举哀说：‘哀哉！我主啊。’这话是我说的。这是耶和华说的。”
JER|34|6|于是， 耶利米 先知在 耶路撒冷 把这一切话告诉 犹大 王 西底家 。
JER|34|7|那时， 巴比伦 王的军队正攻打 耶路撒冷 ，又攻打 犹大 仅存的城镇，就是 拉吉 和 亚西加 ；原来 犹大 的坚固城只剩下这两座。
JER|34|8|西底家 王与 耶路撒冷 的众百姓立约，要他们宣告自由，叫各人释放自己的仆人和婢女，使 希伯来 的男人和女人得自由，谁也不可使他的 犹大 弟兄作奴仆。这事以后，耶和华的话临到 耶利米 。
JER|34|9|
JER|34|10|所有前来立约的领袖和众百姓都顺从，各人释放自己的仆人和婢女，使他们得自由，不再叫他们作奴仆。大家都顺从，将仆婢释放了。
JER|34|11|但后来他们又反悔，叫被释放得自由的仆人婢女回来，强迫他们仍为仆婢。
JER|34|12|因此耶和华的话临到 耶利米 ，说：
JER|34|13|“耶和华－ 以色列 的上帝如此说：我将你们祖先从 埃及 地为奴之家领出时，与他们立约说：
JER|34|14|‘你的一个 希伯来 弟兄若卖给你，服事你六年，到第七年你们各人就要释放他自由出去。’只是你们祖先不听我，不侧耳而听。
JER|34|15|如今你们回转，行我眼中看为正的事，各人向邻舍宣告自由，并且在我面前、在称为我名下的殿中立约。
JER|34|16|你们却反悔，亵渎我的名，各人叫所释放得自由的仆人婢女回来，强迫他们仍为仆婢。
JER|34|17|所以耶和华如此说：你们不听从我，各人不向弟兄邻舍宣告自由。看哪！我要向你们宣告自由，把你们自由地交给刀剑、饥荒、瘟疫，并且使地上万国因你们而惊骇。这是耶和华说的。
JER|34|18|那些违背我约的人，就是不遵守在我面前立约之话的，我要使他们成了那劈成两半的牛犊，使人从切块中经过：
JER|34|19|犹大 的领袖、 耶路撒冷 的领袖、官员、祭司，和从牛犊切块中经过的这地的众百姓，
JER|34|20|我必将他们交在仇敌和寻索其命的人手中；他们的尸首必给空中的飞鸟和地上的走兽作食物。
JER|34|21|我必将 犹大 王 西底家 和他的众领袖交在仇敌和寻索其命的人手中，与那暂时离你们而去的 巴比伦 王军队的手中。
JER|34|22|看哪，我要吩咐他们回到这城，攻打这城，将城攻取，用火焚烧；我也要使 犹大 的城镇变为废墟，无人居住。这是耶和华说的。”
JER|35|1|当 约西亚 的儿子 约雅敬 作 犹大 王的时候，耶和华的话临到 耶利米 ，说：
JER|35|2|“你去见 利甲 族的人，吩咐他们，领他们进入耶和华殿的一个房间，给他们酒喝。”
JER|35|3|我就带 哈巴洗尼雅 的孙子 雅利米雅 的儿子 雅撒尼亚 ，和他的兄弟，并他所有的儿子，以及 利甲 全族的人，
JER|35|4|领他们到耶和华的殿，进入 伊基大利 的儿子神人 哈难 儿子们的房间；那房间靠近官长的房间，在 沙龙 之子门口的守卫 玛西雅 的房间上面。
JER|35|5|于是我在 利甲 族的人面前摆设盛满了酒的碗和杯，对他们说：“请喝酒。”
JER|35|6|他们却说：“我们不喝酒，因为我们祖先 利甲 的儿子 约拿达 曾吩咐我们说：‘你们与你们的子孙永不可喝酒，
JER|35|7|不可盖房子，不可撒种，也不可栽葡萄园，连拥有都不可；但一生的年日要住帐棚，使你们的日子在寄居的地面上得以长久。’
JER|35|8|凡我们祖先 利甲 的儿子 约拿达 所吩咐我们的话，我们都听从了。我们和我们的妻子儿女一生的年日都不喝酒，
JER|35|9|不盖房子居住，我们也没有葡萄园、田地和种子；
JER|35|10|但住在帐棚里，听从并遵行我们祖先 约拿达 所吩咐我们的一切话。
JER|35|11|巴比伦 王 尼布甲尼撒 上来攻打这地的时候，我们说：‘来吧，我们到 耶路撒冷 去，躲避 迦勒底 的军队和 亚兰 的军队。’这样，我们才住在 耶路撒冷 。”
JER|35|12|耶和华的话临到 耶利米 ，说：
JER|35|13|“万军之耶和华－ 以色列 的上帝如此说：你去对 犹大 人和 耶路撒冷 的居民说，你们不肯领受训诲，听从我的话吗？这是耶和华说的。
JER|35|14|利甲 的儿子 约拿达 所吩咐他子孙不可喝酒的话，他们已经遵守了；他们因为听从祖先的吩咐，直到今日都不喝酒。至于我，我一再警戒你们，你们却不肯听从我。
JER|35|15|我一再差遣我的仆人众先知到你们那里去，说：‘你们各人当回头离开恶道，改正行为，不再随从事奉别神，如此，就必住在我所赐给你们和你们祖先的地上。’只是你们不侧耳而听，也不听我。
JER|35|16|利甲 的儿子 约拿达 的子孙能遵守祖先所吩咐他们的命令，这百姓却不肯听从我！
JER|35|17|因此，耶和华－万军之上帝、 以色列 的上帝如此说：看哪，我要使我所说的一切灾祸临到 犹大 人和 耶路撒冷 所有的居民。因为我向他们说话，他们不听从；我呼唤他们，他们也没有回应。”
JER|35|18|耶利米 对 利甲 族的人说：“万军之耶和华－ 以色列 的上帝如此说：因你们听从你们祖先 约拿达 的吩咐，谨守他的一切命令，照他所吩咐的去做，
JER|35|19|所以万军之耶和华－ 以色列 的上帝如此说： 利甲 的儿子 约拿达 必永远不断有人侍立在我面前。”
JER|36|1|约西亚 的儿子 犹大 王 约雅敬 第四年，有这话从耶和华临到 耶利米 ，说：
JER|36|2|“你要取一书卷，把我对你所说攻击 以色列 和 犹大 ，并各国的一切话，从我对你说话的那日，就是从 约西亚 的日子起直到今日，都写在其上；
JER|36|3|或者 犹大 家听见我想要降给他们的一切灾祸，各人就回转离开恶道，我就赦免他们的罪孽和罪恶。”
JER|36|4|耶利米 召了 尼利亚 的儿子 巴录 来； 巴录 就从 耶利米 口中，把耶和华对 耶利米 所说的一切话写在书卷上。
JER|36|5|耶利米 吩咐 巴录 说：“我被禁止，不能进耶和华的殿。
JER|36|6|所以你要趁禁食的日子进入耶和华的殿中，把耶和华的话，就是你从我口中写在书卷上的话，念给百姓和所有从各城镇前来的 犹大 人亲耳听；
JER|36|7|或者他们的恳求达到耶和华面前，各人回转离开恶道，因为耶和华向这百姓所说要发的怒气和愤怒实在很大。”
JER|36|8|尼利亚 的儿子 巴录 就照 耶利米 先知所吩咐的一切去做，在耶和华殿中宣读书卷上耶和华的话。
JER|36|9|约西亚 的儿子 犹大 王 约雅敬 第五年九月， 耶路撒冷 的众百姓和那从 犹大 城镇前来 耶路撒冷 的众百姓，在耶和华面前宣告禁食，
JER|36|10|巴录 就在耶和华殿的上院，靠近耶和华殿的 新门 口， 沙番 的儿子 基玛利雅 文士的房间里，宣读书卷上 耶利米 的话给众百姓亲耳听。
JER|36|11|沙番 的孙子 基玛利雅 的儿子 米该亚 听见书卷上耶和华的一切话，
JER|36|12|就下到王宫，进入书记的房间。看哪，所有的官长都坐在那里，包括 以利沙玛 文士、 示玛雅 的儿子 第莱雅 、 亚革波 的儿子 以利拿单 、 沙番 的儿子 基玛利雅 、 哈拿尼雅 的儿子 西底家 和其余的官长。
JER|36|13|米该亚 向他们述说他所听见的一切话，就是当 巴录 向众百姓宣读那书卷时亲耳听见的。
JER|36|14|官长们就派 犹底 ，就是 古示 的曾孙， 示利米雅 的孙子， 尼探雅 的儿子到 巴录 那里，对他说：“你把你所念给百姓听的书卷拿在手里，到我们这里来。” 尼利亚 的儿子 巴录 就手拿书卷到他们那里来。
JER|36|15|他们对他说：“请坐下，念给我们亲耳听。” 巴录 就念给他们亲耳听。
JER|36|16|他们听见这一切话就害怕，面面相觑，对 巴录 说：“我们必须将这一切话禀告王。”
JER|36|17|他们问 巴录 说：“请你告诉我们，你怎样从他口中写下这一切话呢？”
JER|36|18|巴录 回答说：“他向我口述这一切话，我就用笔墨把它写在书卷上。”
JER|36|19|众官长对 巴录 说：“你和 耶利米 要去躲起来，不可叫人知道你们躲在哪里。”
JER|36|20|众官长把书卷留在 以利沙玛 文士的房间里，然后进院见王，把这一切话说给王听。
JER|36|21|王就派 犹底 去拿这书卷来；他就从 以利沙玛 文士的房间内取来，念给王和侍立在王左右的众官长亲耳听。
JER|36|22|那时正是九月，王坐在过冬的房屋里，王前面有燃烧的火盆 。
JER|36|23|犹底 念了三、四段 ，王就用文士的刀把书卷割破，丢在火盆里，直到全卷在火中烧尽了。
JER|36|24|王和听见这一切话的臣仆都不惧怕，也不撕裂衣服。
JER|36|25|以利拿单 和 第莱雅 ，并 基玛利雅 恳求王不要烧这书卷，王却不听。
JER|36|26|王吩咐王 的儿子 耶拉篾 、 亚斯列 的儿子 西莱雅 和 亚伯叠 的儿子 示利米雅 ，去捉拿 巴录 文士和 耶利米 先知；耶和华却将他们隐藏起来。
JER|36|27|王烧了有 巴录 从 耶利米 口中所写之话的书卷以后，耶和华的话临到 耶利米 ，说：
JER|36|28|“你再取一书卷，将 犹大 王 约雅敬 所烧前一卷书上原有的一切话写在上面。
JER|36|29|论到 犹大 王 约雅敬 你要说，耶和华如此说：你烧了这书卷，说：‘你为什么在上面写着， 巴比伦 王必要来毁灭这地，使这地绝了人民和牲畜呢？’
JER|36|30|所以耶和华论到 犹大 王 约雅敬 说：他后裔中必没有人坐在 大卫 的宝座上；他的尸首必被抛弃，白天受炎热，黑夜受寒霜。
JER|36|31|我必因他和他后裔，并他臣仆的罪孽惩罚他们。我要使我所说的一切灾祸临到他们和 耶路撒冷 的居民，并 犹大 人；只是他们不肯听从。”
JER|36|32|于是， 耶利米 又取一书卷交给 尼利亚 的儿子 巴录 文士，他就从 耶利米 的口中写了 犹大 王 约雅敬 在火中所烧书卷上的一切话，另外又添了许多相仿的话。
JER|37|1|约西亚 的儿子 西底家 接续 约雅敬 的儿子 哥尼雅 作王，因为 巴比伦 王 尼布甲尼撒 立他在 犹大 地作王。
JER|37|2|但 西底家 、他的臣仆和这地的百姓都不听从耶和华藉 耶利米 先知所说的话。
JER|37|3|西底家 王派 示利米雅 的儿子 犹甲 和 玛西雅 的儿子 西番雅 祭司，去见 耶利米 先知，说：“求你为我们祈求耶和华－我们的上帝。”
JER|37|4|那时 耶利米 仍在百姓中进出，因为他们还没有把他囚在监里。
JER|37|5|法老的军队已经从 埃及 出来，那围困 耶路撒冷 的 迦勒底 人听见这风声，就拔营离开 耶路撒冷 去了。
JER|37|6|耶和华的话临到 耶利米 先知，说：
JER|37|7|“耶和华－ 以色列 的上帝如此说：你们要对派你们来求问我的 犹大 王如此说：‘看哪，那出来帮助你们的法老军队必回 埃及 本国去。
JER|37|8|迦勒底 人必再来攻打这城，并要攻下，用火焚烧。
JER|37|9|耶和华如此说：你们不要自欺说“ 迦勒底 人必定离开我们”，因为他们必不离开。
JER|37|10|你们即使击败与你们争战的 迦勒底 全军，他们当中剩下受伤的人也必各自从帐棚里起来，用火焚烧这城。’”
JER|37|11|迦勒底 的军队因躲避法老的军队，拔营离开 耶路撒冷 的时候，
JER|37|12|耶利米 离开 耶路撒冷 ，往 便雅悯 地去，要在那里从百姓当中取得自己的地产。
JER|37|13|他到了 便雅悯门 ，那里的守门官名叫 伊利雅 ，是 哈拿尼亚 的孙子， 示利米雅 的儿子，他逮捕 耶利米 先知，说：“你是去投降 迦勒底 人的！”
JER|37|14|耶利米 说：“你这是谎话，我并不是去投降 迦勒底 人。” 伊利雅 不听 耶利米 的话，就逮捕他，把他带到官长那里。
JER|37|15|官长们恼怒 耶利米 ，打了他，把他囚在 约拿单 文士的房屋中，因为他们把这屋子当作监牢。
JER|37|16|耶利米 来到地牢，进入牢房，在那里拘留多日。
JER|37|17|西底家 王差人提他出来，在自己的宫内私下问他说：“有什么话从耶和华临到没有？” 耶利米 说：“有！”又说：“你必被交在 巴比伦 王手中。”
JER|37|18|耶利米 又对 西底家 王说：“我在什么事上得罪你，或你的臣仆，或这百姓，你们竟将我囚在监里呢？
JER|37|19|对你们预言‘ 巴比伦 王必不来攻击你们和这地’的先知在哪里呢？
JER|37|20|主－我的王啊，现在求你垂听，允准我在你面前的恳求：不要把我送回 约拿单 文士的房屋中，免得我死在那里。”
JER|37|21|于是 西底家 王下令，他们就把 耶利米 交在护卫兵的院中，每天从饼店街取一个饼给他，直到城中所有的饼都用尽了。这样， 耶利米 仍拘留在护卫兵的院中。
JER|38|1|玛坦 的儿子 示法提雅 、 巴施户珥 的儿子 基大利 、 示利米雅 的儿子 犹甲 、 玛基雅 的儿子 巴示户珥 听见 耶利米 对众百姓所说的话，说：
JER|38|2|“耶和华如此说：留在这城里的必遭刀剑、饥荒、瘟疫而死，但归向 迦勒底 人的必得存活；至少能保全自己的性命，得以存活。
JER|38|3|耶和华如此说：这城必要交在 巴比伦 王军队的手中，他必攻下这城。”
JER|38|4|于是官长们对王说：“求你把这人处死，因他向城里剩下的士兵和众人说这样的话，使他们的手发软。这人不是为这百姓求平安，而是叫他们受灾祸。”
JER|38|5|西底家 王说：“看哪，他在你们手中，王不能反对你们所做的事。”
JER|38|6|他们就拿住 耶利米 ，把他丢在王 的儿子 玛基雅 的井里；那口井在护卫兵的院中。他们用绳子把 耶利米 缒下去，井里没有水，只有淤泥， 耶利米 就陷在淤泥中。
JER|38|7|在王宫里的太监 古实 人 以伯．米勒 ，听见他们把 耶利米 丢进井里，那时王坐在 便雅悯门 前。
JER|38|8|以伯．米勒 从王宫里出来，对王说：
JER|38|9|“主－我的王啊，这些人向 耶利米 先知一味地行恶，把他丢在井里；他在那里必因饥饿而死，因为城里不再有粮食了。”
JER|38|10|王就吩咐 古实 人 以伯．米勒 说：“你从这里带领三十人，趁 耶利米 先知还没死，把他从井里拉上来。”
JER|38|11|于是 以伯．米勒 带领这些人同去，进入王宫，到库房以下 ，从那里取了些碎布和破衣服，用绳子缒下去，到井里 耶利米 那里。
JER|38|12|古实 人 以伯．米勒 对 耶利米 说：“你用这些碎布和破衣服放在绳子上，垫你的腋下。” 耶利米 就照样做。
JER|38|13|这样，他们用绳子将 耶利米 从井里拉上来。 耶利米 仍在护卫兵的院中。
JER|38|14|西底家 王差人将 耶利米 先知带进耶和华殿的第三个门，到王那里去。王对 耶利米 说：“我要问你一件事，你一点都不可向我隐瞒。”
JER|38|15|耶利米 对 西底家 说：“我若告诉你，你岂不是一定要把我处死吗？我若劝你，你必不听我。”
JER|38|16|西底家 王就私下对 耶利米 说：“我指着那造我们生命之永生的耶和华起誓：我必不把你处死，也不将你交在寻索你命的人手中。”
JER|38|17|耶利米 对 西底家 说：“耶和华－万军之上帝、 以色列 的上帝如此说：你若归顺 巴比伦 王的官长，你的命就必存活，这城也不致被火焚烧，你和你的全家都必存活。
JER|38|18|你若不归顺 巴比伦 王的官长，这城必交在 迦勒底 人手中。他们必用火焚烧，你也不得脱离他们的手。”
JER|38|19|西底家 王对 耶利米 说：“我怕那些投降 迦勒底 人的 犹大 人，恐怕 迦勒底 人把我交在他们手中，他们就戏弄我。”
JER|38|20|耶利米 说：“ 迦勒底 人必不把你交出。求你听从我对你所说耶和华的话，这样对你有好处，你的命也必存活。
JER|38|21|你若不肯归顺，耶和华指示我的话是这样：
JER|38|22|看哪， 犹大 王宫里所留下来的妇女必被带到 巴比伦 王的官长那里。这些妇女要说： 你知己的朋友引诱你， 他们胜过你； 你的脚陷入淤泥， 他们却离弃你。
JER|38|23|“人必将你的后妃和你的儿女带到 迦勒底 人那里；你也不得脱离他们的手，必被 巴比伦 王的手捉住，这城也必被火焚烧 。”
JER|38|24|西底家 对 耶利米 说：“不要让人知道这些对话，你就不至于死。
JER|38|25|官长们若听见我跟你说话，到你那里对你说：‘告诉我们，你对王说了什么话，王又向你说了什么；不可向我们隐瞒，否则我们就要杀你。’
JER|38|26|你就对他们说：‘我在王面前恳求不要把我送回 约拿单 的房屋，免得我死在那里。’”
JER|38|27|随后官长们到 耶利米 那里，问他，他就照王所吩咐的一切话回答他们。他们就不再问他，因为事情没有泄漏。
JER|38|28|于是 耶利米 仍在护卫兵的院中，直到 耶路撒冷 被攻下的日子。当 耶路撒冷 被攻下时，他仍在那里。
JER|39|1|犹大 王 西底家 第九年十月， 巴比伦 王 尼布甲尼撒 率领全军前来围困 耶路撒冷 。
JER|39|2|西底家 十一年四月初九日，城被攻破。
JER|39|3|耶路撒冷 被攻下的时候， 巴比伦 王的众官长， 尼甲．沙利薛 、 三甲．尼波 、 撒西金 将军 、 尼甲．沙利薛 将军 ，并 巴比伦 王其余的官长都来坐在 中门 。
JER|39|4|犹大 王 西底家 和所有士兵看见他们，就在夜间从靠近王的花园、两城墙中间的门逃跑出城，往 亚拉巴 逃去。
JER|39|5|迦勒底 的军队追赶他们，在 耶利哥 的平原追上 西底家 ，将他逮住，带到 哈马 地的 利比拉 、 巴比伦 王 尼布甲尼撒 那里； 尼布甲尼撒 就判他的罪。
JER|39|6|在 利比拉 ， 巴比伦 王在 西底家 眼前杀了他的儿女； 巴比伦 王又杀了 犹大 所有的贵族，
JER|39|7|并且挖了 西底家 的眼睛，用铜链锁住他，要带到 巴比伦 去。
JER|39|8|迦勒底 人用火焚烧王宫和百姓的房屋，又拆毁 耶路撒冷 的城墙。
JER|39|9|那时， 尼布撒拉旦 护卫长把城里所剩下的百姓和投降他的降民，以及其余的百姓都掳到 巴比伦 去了。
JER|39|10|尼布撒拉旦 护卫长却把百姓中一无所有的穷人留在 犹大 地，当时就赏给他们葡萄园和田地 。
JER|39|11|巴比伦 王 尼布甲尼撒 为了 耶利米 ，嘱咐 尼布撒拉旦 护卫长：
JER|39|12|“你领他去，好好地看待他，切不可害他；他对你怎么说，你就向他怎样做。”
JER|39|13|尼布撒拉旦 护卫长和 尼布沙斯班 将军 、 尼甲．沙利薛 将军 ，并 巴比伦 王众官长，
JER|39|14|派人把 耶利米 从护卫兵的院中提出来，交给 沙番 的孙子， 亚希甘 的儿子 基大利 ，让他自由进出屋子；于是 耶利米 住在百姓中间。
JER|39|15|耶利米 还囚在护卫兵院中的时候，耶和华的话临到他，说：
JER|39|16|“你去告诉 古实 人 以伯．米勒 说，万军之耶和华－ 以色列 的上帝如此说：看哪，我说降祸不降福的话必临到这城，到那时必在你面前实现。
JER|39|17|到那日我必拯救你，你必不致交在你所怕的人手中。这是耶和华说的。
JER|39|18|我定要搭救你，你必不致倒在刀下，却要保全自己的性命，因你倚靠我。这是耶和华说的。”
JER|40|1|耶利米 被链子锁在 耶路撒冷 和 犹大 被掳到 巴比伦 的人中， 尼布撒拉旦 护卫长把他从 拉玛 提出来，释放他以后，耶和华的话临到 耶利米 。
JER|40|2|护卫长提 耶利米 来，对他说：“耶和华－你的上帝曾说要降这灾祸给此地。
JER|40|3|耶和华照他所说的做了，已使这灾祸临到；因你们得罪耶和华，不听从他的话，所以这事临到你们。
JER|40|4|看哪，现在我解开你手上的链子，你若看与我同往 巴比伦 去好，就可以去，我必厚待你；你若看与我同往 巴比伦 去不好，就不必去。看哪，全地在你面前，你以为哪里美好，哪里合宜，只管去吧
JER|40|5|─ 耶利米 尚未回去 ─你可以回到 巴比伦 王所立管理 犹大 城镇的 沙番 的孙子， 亚希甘 的儿子 基大利 那里去，在他那里住在百姓当中。不然，你看哪里合宜就可以去。”于是护卫长送他粮食和礼物，释放了他。
JER|40|6|耶利米 就来到 米斯巴 ， 亚希甘 的儿子 基大利 那里去，与他同住，住在留于境内的百姓当中。
JER|40|7|在乡间所有的军官和属他们的人，听见 巴比伦 王立了 亚希甘 的儿子 基大利 作当地的省长，并将没有掳到 巴比伦 的男人、妇女、孩童和当地极穷的人全交给他，
JER|40|8|于是 尼探雅 的儿子 以实玛利 ， 加利亚 的两个儿子 约哈难 和 约拿单 ， 单户篾 的儿子 西莱雅 ，并 尼陀法 人 以斐 的众子， 玛迦 人的儿子 耶撒尼亚 ，和属他们的人，都来到 米斯巴 的 基大利 那里。
JER|40|9|沙番 的孙子， 亚希甘 的儿子 基大利 向他们和属他们的人起誓说：“不要怕服事 迦勒底 人，只管住在这地，服事 巴比伦 王，就可以得福。
JER|40|10|至于我，我要住在 米斯巴 ，侍候那些到我们这里来的 迦勒底 人；只是你们当积蓄酒、油和夏天的果子，收藏在器皿里，并住在你们所占的城镇中。”
JER|40|11|在 摩押 地和 亚扪 人当中，在 以东 地和各国，所有的 犹大 人听见 巴比伦 王留下一些 犹大 人，并立 沙番 的孙子、 亚希甘 的儿子 基大利 管理他们，
JER|40|12|所有的 犹大 人就从被赶到的各处回来，到 犹大 地 米斯巴 的 基大利 那里。他们积蓄了许多的酒，并夏天的果子。
JER|40|13|加利亚 的儿子 约哈难 和在乡间的军官来到 米斯巴 的 基大利 那里，
JER|40|14|对他说：“ 亚扪 人的王 巴利斯 派 尼探雅 的儿子 以实玛利 来谋害你的命，你知道吗？” 亚希甘 的儿子 基大利 却不相信他们的话。
JER|40|15|加利亚 的儿子 约哈难 在 米斯巴 私下对 基大利 说：“求你容我去杀 尼探雅 的儿子 以实玛利 ，必无人知道。何必让他害你的命，使聚集到你这里来的 犹大 人都分散，以致 犹大 剩余的人都灭亡呢？”
JER|40|16|亚希甘 的儿子 基大利 对 加利亚 的儿子 约哈难 说：“你不可做这事，你所论 以实玛利 的话是假的。”
JER|41|1|七月中，王的大臣，就是王室后裔 以利沙玛 的孙子、 尼探雅 的儿子 以实玛利 带着十个人，来到 米斯巴 ， 亚希甘 的儿子 基大利 那里；他们在 米斯巴 一同吃饭。
JER|41|2|尼探雅 的儿子 以实玛利 和同他来的那十个人起来，用刀击杀 沙番 的孙子， 亚希甘 的儿子 基大利 ，就是 巴比伦 王所立为当地省长的，把他杀死。
JER|41|3|以实玛利 把所有在 米斯巴 与 基大利 一起的 犹大 人，以及他们在那里所遇见的 迦勒底 人和士兵都杀了。
JER|41|4|他杀了 基大利 的第二天，还没有人知道的时候，
JER|41|5|有八十人从 示剑 、 示罗 和 撒玛利亚 前来，胡须剃去，衣服撕裂，身体划破，手拿素祭和乳香，要奉到耶和华的殿。
JER|41|6|尼探雅 的儿子 以实玛利 从 米斯巴 出来迎接他们，随走随哭，遇见了他们，就对他们说：“你们可以到 亚希甘 的儿子 基大利 那里。”
JER|41|7|他们到了城中， 尼探雅 的儿子 以实玛利 和与他一起的人就把他们杀了，丢在坑里。
JER|41|8|只是他们中间有十个人对 以实玛利 说：“不要杀我们，因为我们有许多大麦、小麦、油和蜜藏在田间。”于是他住手，没有在弟兄中间杀他们。
JER|41|9|以实玛利 把那些因 基大利 事件所杀之人的尸首都丢在坑里；这坑是从前 亚撒 王因怕 以色列 王 巴沙 所挖的。 尼探雅 的儿子 以实玛利 把那些被杀的人填满了坑。
JER|41|10|以实玛利 把 米斯巴 剩下的人，就是众公主和仍住在 米斯巴 所有的百姓都掳去，他们原是 尼布撒拉旦 护卫长交给 亚希甘 的儿子 基大利 的。 尼探雅 的儿子 以实玛利 掳了他们，要到 亚扪 人那里去。
JER|41|11|加利亚 的儿子 约哈难 和与他一起的军官，听见 尼探雅 的儿子 以实玛利 所做的一切恶事，
JER|41|12|就带领众人前往，要和 尼探雅 的儿子 以实玛利 争战，他们在 基遍 的大水池 旁遇见他。
JER|41|13|在 以实玛利 那里的众人看见 加利亚 的儿子 约哈难 和与他一起的军官，就都欢喜。
JER|41|14|这样， 以实玛利 从 米斯巴 所掳去的众人都转而归向 加利亚 的儿子 约哈难 。
JER|41|15|尼探雅 的儿子 以实玛利 和八个人脱离 约哈难 的手，逃到 亚扪 人那里去。
JER|41|16|尼探雅 的儿子 以实玛利 杀了 亚希甘 的儿子 基大利 ，从 米斯巴 把所有幸存的百姓、士兵、妇女、孩童、太监掳到 基遍 之后， 加利亚 的儿子 约哈难 和与他一起的军官把他们都抢回来，
JER|41|17|带到靠近 伯利恒 的 基罗特金罕 住下，要到 埃及 去，
JER|41|18|躲避 迦勒底 人。他们惧怕 迦勒底 人，因为 尼探雅 的儿子 以实玛利 杀了 巴比伦 王所立管理那地的 亚希甘 的儿子 基大利 。
JER|42|1|众军官和 加利亚 的儿子 约哈难 ，并 何沙雅 的儿子 耶撒尼亚 以及众百姓，从最小的到最大的都进前来，
JER|42|2|对 耶利米 先知说：“请你准我们在你面前祈求，为我们这幸存的人向耶和华－你的上帝祷告。我们本来众多，现在剩下的极少，这是你亲眼看见的。
JER|42|3|愿耶和华－你的上帝指示我们当走的路，当做的事。”
JER|42|4|耶利米 先知对他们说：“我已经听见了，看哪，我必照你们的话向耶和华－你们的上帝祷告。耶和华无论回答什么，我都必告诉你们，绝不隐瞒。”
JER|42|5|于是他们对 耶利米 说：“我们若不照耶和华－你上帝差遣你说的一切话去做，愿耶和华在我们中间作真实可靠的见证。
JER|42|6|我们请你到耶和华－我们的上帝面前，他说的无论是好是歹，我们都必听从；因为我们听从耶和华－我们上帝的话，就可以得福。”
JER|42|7|过了十天，耶和华的话临到 耶利米 。
JER|42|8|他就将 加利亚 的儿子 约哈难 和与他一起所有的军官和百姓，从最小的到最大的都召来，
JER|42|9|对他们说：“你们请我到耶和华－ 以色列 的上帝面前为你们祈求，他如此说：
JER|42|10|‘你们若仍留在这地，我就建立你们，必不拆毁；栽植你们，必不拔出；因我为所降与你们的灾祸感到遗憾。
JER|42|11|不要怕你们所惧怕的 巴比伦 王。不要怕他！因为我与你们同在，要拯救你们脱离他的手。这是耶和华说的。
JER|42|12|我要向你们施怜悯，他 就怜悯你们，使你们归回本地。’
JER|42|13|倘若你们说：‘我们不留在这地’，不听从耶和华－你们上帝的话，
JER|42|14|说：‘我们不留在这地，却要进入 埃及 地，在那里我们看不见战争，听不见角声，也不致缺食挨饿；我们要住在那里。’
JER|42|15|幸存的 犹大 人哪，你们现在要听耶和华的话；万军之耶和华－ 以色列 的上帝如此说：‘你们若定意进入 埃及 ，在那里寄居，
JER|42|16|你们所惧怕的刀剑在 埃及 地必追上你们，你们所惧怕的饥荒在 埃及 要紧紧跟随你们，你们必死在那里。
JER|42|17|凡定意进入 埃及 在那里寄居的，必遭刀剑、饥荒、瘟疫而死，无一人存留，得以逃脱我所降与他们的灾祸。’
JER|42|18|“万军之耶和华－ 以色列 的上帝如此说：‘我怎样将我的怒气和愤怒倾倒在 耶路撒冷 的居民身上，你们进入 埃及 的时候，我也必照样将我的愤怒倾倒在你们身上，以致你们受辱骂、惊骇、诅咒、羞辱，并且不得再看见这地方。’
JER|42|19|幸存的 犹大 人哪，耶和华论到你们说：‘不要进入 埃及 。’你们要确实知道，我今日已警戒你们了。
JER|42|20|你们行诡诈害自己；因为你们请我到耶和华－你们上帝那里，说：‘请你为我们向耶和华－我们的上帝祷告，你把耶和华－我们上帝所说的一切告诉我们，我们就必遵行。’
JER|42|21|我今日把这话告诉你们，你们却不听耶和华－你们上帝为这一切事差我到你们那里所说的话。
JER|42|22|现在你们要确实知道，你们在所要去的寄居之地必遭刀剑、饥荒、瘟疫而死。”
JER|43|1|耶利米 向众百姓说完了耶和华－他们上帝一切的话，就是耶和华－他们上帝差他去说的这一切话，
JER|43|2|何沙雅 的儿子 亚撒利雅 和 加利亚 的儿子 约哈难 ，以及所有狂傲的人，就对 耶利米 说：“你说谎！耶和华－我们的上帝并没有差遣你说：‘你们不可进入 埃及 ，在那里寄居。’
JER|43|3|这是 尼利亚 的儿子 巴录 挑唆你害我们，要把我们交在 迦勒底 人手中，使我们被杀或被掳到 巴比伦 去。”
JER|43|4|加利亚 的儿子 约哈难 和所有的军官、百姓，都不肯听从耶和华的话留在 犹大 地。
JER|43|5|加利亚 的儿子 约哈难 和所有的军官却将幸存的 犹大 人，就是从被赶到的各国回来，在 犹大 地寄居的男人、妇女、孩童和众公主，并 尼布撒拉旦 护卫长留在 沙番 的孙子， 亚希甘 的儿子 基大利 那里的众人，与 耶利米 先知，以及 尼利亚 的儿子 巴录 ，
JER|43|6|
JER|43|7|都带入 埃及 地，到了 答比匿 ；这是因他们不肯听从耶和华的话。
JER|43|8|在 答比匿 ，耶和华的话临到 耶利米 ，说：
JER|43|9|“你要在 犹大 人眼前用手拿几块大石头，藏在 答比匿 法老的宫门砌砖的石墩上，
JER|43|10|对他们说：‘万军之耶和华－ 以色列 的上帝如此说：看哪，我必召我的仆人 巴比伦 王 尼布甲尼撒 前来，安置他的宝座在所藏的这些石头上；他要在其上支搭华丽的帐幕。
JER|43|11|他要来攻击 埃及 地： 定为死亡的，必致死亡； 定为掳掠的，必遭掳掠； 定为刀杀的，必被刀杀。
JER|43|12|我要用火点燃 埃及 众神明的庙宇， 巴比伦 王要焚烧庙宇，掳去神像；他要围住 埃及 地，好像牧人披上外衣，从那里安然而去。
JER|43|13|他必打碎 埃及 地 伯．示麦 的柱像，用火焚烧 埃及 众神明的庙宇。’”
JER|44|1|有话临到 耶利米 ，论到住 埃及 地所有的 犹大 人，就是住在 密夺 、 答比匿 、 挪弗 、 巴特罗 境内的 犹大 人，说：
JER|44|2|“万军之耶和华－ 以色列 的上帝如此说：我所降与 耶路撒冷 和 犹大 各城的一切灾祸，你们都看见了。看哪，那些城镇今日荒凉，无人居住；
JER|44|3|这是因居民所行的恶，去烧香事奉别神，就是他们和你们，以及你们列祖所不认识的神明，惹我发怒。
JER|44|4|我一再差遣我的仆人众先知去，说：你们切不可行我所厌恶这可憎之事。
JER|44|5|他们却不听从，不侧耳而听，也不转离恶事，仍向别神烧香。
JER|44|6|因此，我的怒气和愤怒都倾倒出来，在 犹大 城镇和 耶路撒冷 街市上燃起，以致它们都荒废凄凉，正如今日一样。
JER|44|7|现在耶和华－万军之上帝、 以色列 的上帝如此说：你们为何做这大恶自害己命，使你们的男人、妇女、孩童和吃奶的都从 犹大 剪除，不留一人呢？
JER|44|8|你们以手所做的，在寄居的 埃及 地向别神烧香，惹我发怒，使你们被剪除，在天下万国中受诅咒羞辱。
JER|44|9|你们祖先的恶行， 犹大 诸王和后妃的恶行，你们自己和你们妻子的恶行，就是在 犹大 地和 耶路撒冷 街市上所做的，你们都忘了吗？
JER|44|10|到如今你们还不懊悔，不惧怕，不肯遵行我在你们和你们祖先面前所设立的法度律例。
JER|44|11|“所以万军之耶和华－ 以色列 的上帝如此说：看哪，我必向你们变脸降灾，剪除 犹大 众人。
JER|44|12|我必使那定意进入 埃及 地、在那里寄居的，就是幸存的 犹大 人，尽都灭绝。他们必在 埃及 地仆倒，因刀剑饥荒灭绝，从最小的到最大的都必遭刀剑饥荒而死，甚至受辱骂、惊骇、诅咒、羞辱。
JER|44|13|我怎样用刀剑、饥荒、瘟疫惩罚 耶路撒冷 ，也必照样惩罚那些住在 埃及 地的 犹大 人。
JER|44|14|那进入 埃及 地、在那里寄居的，就是幸存的 犹大 人，都不得逃脱，也不得归回 犹大 地。他们心中很想归回，居住在那里；但除了少数逃脱的以外，都不得归回。”
JER|44|15|那些知道自己妻子向别神烧香的男人，与站在那里的一大群妇女，就是住 埃及 地 巴特罗 所有的百姓，回答 耶利米 说：
JER|44|16|“论到你奉耶和华的名向我们所说的话，我们必不听从。
JER|44|17|我们定要照我们口中所说的一切话去做，向天后烧香，献浇酒祭，按着我们与我们祖先、君王、官长在 犹大 城镇和 耶路撒冷 街市上素常所做的一样；因为那时我们得以吃饱、享福乐，并未遇见灾祸。
JER|44|18|自从我们停止向天后烧香，献浇酒祭，我们倒缺乏这一切，又因刀剑饥荒灭绝。”
JER|44|19|妇女们说 ：“我们向天后烧香，献浇酒祭，做天后像的饼供奉它，向它献浇酒祭，难道我们的丈夫没有参与吗？”
JER|44|20|耶利米 对这样回答他的男人和妇女说：
JER|44|21|“你们与你们祖先、君王、官长，以及这地的百姓，在 犹大 城镇和 耶路撒冷 街市上所烧的香，耶和华岂不记得，放在他心上吗？
JER|44|22|耶和华因你们所行的恶、所做可憎的事，不能再容忍，所以使你们的地荒凉，受惊骇诅咒，无人居住，正如今日一样。
JER|44|23|你们烧香，得罪耶和华，不听耶和华的话，不遵行他的律法、条例、法度，所以你们遭遇这灾祸，正如今日一样。”
JER|44|24|耶利米 又对众百姓和妇女说：“所有在 埃及 地的 犹大 人哪，当听耶和华的话。
JER|44|25|万军之耶和华－ 以色列 的上帝如此说：你们和你们的妻子口中说过、手里做到，说：‘我们定要向天后还愿，向它烧香，献浇酒祭。’现在你们尽管坚定所许的愿，去还愿吧！
JER|44|26|所有住 埃及 地的 犹大 人哪，当听耶和华的话。耶和华说：看哪，我指着我至大的名起誓，在 埃及 全地，我的名必不再被 犹大 任何人的口呼喊：‘我指着主－永生的耶和华起誓。’
JER|44|27|看哪，我看守他们，为要降祸不降福；在 埃及 地的 犹大 人必因刀剑、饥荒而灭亡，直到灭绝。
JER|44|28|从 埃及 地能脱离刀剑、归回 犹大 地的人数很少。那进入 埃及 地、在那里寄居的，就是幸存的 犹大 人，必知道是谁的话站得住，是我的话呢，还是他们的话。
JER|44|29|我在这地方惩罚你们，必有预兆，使你们知道我降祸给你们的话必站得住。这是耶和华说的。
JER|44|30|耶和华如此说：看哪，我必将 埃及 王 合弗拉 法老交在他仇敌和寻索其命的人手中，像我将 犹大 王 西底家 交在他仇敌和寻索其命的 巴比伦 王 尼布甲尼撒 手中一样。”
JER|45|1|约西亚 的儿子 犹大 王 约雅敬 第四年， 尼利亚 的儿子 巴录 把 耶利米 先知口中所说的话写在书上； 耶利米 对 巴录 说：
JER|45|2|“ 巴录 啊，耶和华－ 以色列 的上帝说：
JER|45|3|你曾说：‘哀哉！耶和华使我愁上加愁，我因呻吟而困乏，不得安歇。’
JER|45|4|你要这样告诉他，耶和华如此说：看哪，我所建立的，我必拆毁；我所栽植的，我必拔出；在全地我都如此行。
JER|45|5|你为自己图谋大事吗？不要图谋！看哪，我必使灾祸临到凡有血肉之躯的。但你无论往哪里去，我要保全你的性命。这是耶和华说的。”
JER|46|1|耶和华论列国的话临到 耶利米 先知。
JER|46|2|论到 埃及 ，关于 埃及 王 尼哥 法老的军队，这军队安营在 幼发拉底河 边的 迦基米施 ，是 巴比伦 王 尼布甲尼撒 在 约西亚 的儿子 犹大 王 约雅敬 第四年所打败的。
JER|46|3|你们要预备大小盾牌， 往前上阵，
JER|46|4|套上车， 骑上马！ 顶盔站立， 磨枪披甲！
JER|46|5|我为何看见他们惊惶， 转身退后呢？ 他们的勇士打败仗， 急忙逃跑，并不回头； 四围都有惊吓！ 这是耶和华说的。
JER|46|6|不要容快跑的逃避， 也不要容勇士逃脱 ； 在北方 幼发拉底河 边， 他们绊跌仆倒。
JER|46|7|这是谁，像 尼罗河 涨溢， 如江河的水翻腾呢？
JER|46|8|埃及 像 尼罗河 涨溢， 如江河的水翻腾。 它说：“我要涨溢遮盖全地； 我要毁灭城镇和其中的居民。
JER|46|9|马匹啊，上去吧！ 战车啊，要疾行！ 手拿盾牌的 古实 和 弗 的勇士， 擅长拉弓的 路德 人，前进吧！”
JER|46|10|那日是万军之主耶和华报仇的日子， 要向敌人报仇。 刀剑必吞吃饱足， 饮血满足； 因为在北方 幼发拉底河 边， 有祭物献给万军之主耶和华。
JER|46|11|少女 埃及 啊， 要上 基列 去取乳香； 你虽服用许多药， 还是徒然，不得治好。
JER|46|12|列国听见你的羞辱， 遍地满了你的哀声； 勇士与勇士彼此相撞， 二人一起跌倒。
JER|46|13|以下是耶和华对 耶利米 先知说的话，论到 巴比伦 王 尼布甲尼撒 要来攻击 埃及 地。
JER|46|14|你们要在 埃及 传扬，在 密夺 报告， 在 挪弗 、 答比匿 宣告说： “要摆好阵势，预备作战， 因为刀剑在你四围施行吞灭。”
JER|46|15|你的壮士为何被扫除呢？ 他们站立不住， 因为耶和华驱逐他们；
JER|46|16|他使多人绊跌，彼此撞倒。 他们说：“起来，让我们回到自己的同胞、 回到自己的出生地去， 好躲避欺压的刀剑。”
JER|46|17|他们在那里称 埃及 王法老 为 “错失良机的夸大者”。
JER|46|18|名为万军之耶和华的君王说： 我指着我的永生起誓： “ 尼布甲尼撒 来的时候， 必像众山之中的 他泊 ， 像海边的 迦密 。”
JER|46|19|住在 埃及 的啊， 要预备被掳时需用的物品； 因为 挪弗 必成为废墟， 被烧毁，无人居住。
JER|46|20|埃及 是肥美的母牛犊； 但来自北方的牛虻来到了！来到了！
JER|46|21|它的佣兵好像圈里的肥牛犊， 他们转身退后， 一齐逃跑，站立不住； 因为他们遭难的日子、 受罚的时刻已经来临。
JER|46|22|它的声音好像蛇在滑行。 敌人要成队而来，如砍伐树木的人， 手拿斧头攻击它。
JER|46|23|虽然它的树林不易穿过， 敌人却要砍伐， 因敌人比蝗虫还多，不可胜数。 这是耶和华说的。
JER|46|24|埃及 必然蒙羞， 被交在北方人的手中。
JER|46|25|万军之耶和华－ 以色列 的上帝说：“看哪，我要惩罚 挪 的 亚扪 和法老、 埃及 和它的神明，以及君王，也要惩罚法老和倚靠他的人。
JER|46|26|我要将他们交给寻索其命之人的手和 巴比伦 王 尼布甲尼撒 与他臣仆的手。但 埃及 日后必再有人居住，与从前一样。这是耶和华说的。”
JER|46|27|我的仆人 雅各 啊，不要惧怕！ 以色列 啊，不要惊惶！ 因我要从远方拯救你， 从被掳之地拯救你的后裔。 雅各 必回来，得享平静安逸， 无人令他害怕。
JER|46|28|我的仆人 雅各 啊，不要惧怕！ 因我与你同在。 我要将那些国灭绝净尽， 就是我赶你去的那些国； 却不将你灭绝净尽， 倒要从宽惩治你， 但绝不能不罚你。 这是耶和华说的。
JER|47|1|在法老攻击 迦萨 之前，耶和华论 非利士 人的话临到 耶利米 先知。
JER|47|2|耶和华如此说： 看哪，有水从北方涨起，成为涨溢的河， 要淹没全地和其中所充满的， 淹没城和城里的居民。 人必呼喊， 境内的居民都必哀号。
JER|47|3|一听见敌人壮马蹄踏的响声、 战车隆隆、车轮轰轰， 为父的手就发软， 不能回头看顾儿女。
JER|47|4|因为日子将到， 耶和华必毁灭所有 非利士 人， 剪除 推罗 、 西顿 仅存的帮助者； 他要毁灭 非利士 人、 迦斐托 海岛剩余的人。
JER|47|5|迦萨 成了光秃， 亚实基伦 归于无有。 平原 中所剩的啊， 你割划自己，要到几时呢？
JER|47|6|耶和华的刀剑哪，你要到几时才止息呢？ 要入鞘，安静不动。
JER|47|7|耶和华吩咐它攻击 亚实基伦 和海边之地， 既已派定它，你 怎能静止不动呢？
JER|48|1|论 摩押 。 万军之耶和华－ 以色列 的上帝如此说： 祸哉， 尼波 ！它要变为废墟。 基列亭 蒙羞被攻取， 米斯迦 蒙羞被毁坏，
JER|48|2|摩押 不再被称赞。 有人在 希实本 设计谋害它： “来吧！我们将它剪除，使它不再成国。” 玛得缅 哪，你也必静默无声； 刀剑必追赶你。
JER|48|3|从 何罗念 有哀号声： “荒凉！大毁灭！”
JER|48|4|“ 摩押 毁灭了！” 它的孩童哀号，使人听见。
JER|48|5|人上 鲁希坡 随走随哭， 因为在 何罗念 的下坡听见毁灭的哀声。
JER|48|6|你们要奔逃，自救己命， 使你们的性命如旷野里的矮树 。
JER|48|7|你因倚靠自己所做的 和自己的财宝，必被攻取。 基抹 和属它的祭司、官长也要一同被掳去。
JER|48|8|那行毁灭的要来到各城， 并无一城幸免。 山谷必败落， 平原必毁坏， 正如耶和华所说的。
JER|48|9|你们要将翅膀给 摩押 ， 使它可以飞去 。 它的城镇必荒凉， 无人居住。
JER|48|10|懒惰不肯为耶和华做事的，必受诅咒；禁止刀剑不见血的，必受诅咒。
JER|48|11|摩押 自幼年以来常享安逸， 如沉淀未被搅动的酒 ， 没有从这器皿倒在那器皿， 也未曾被掳掠过。 因此，它的原味尚存， 香气未变。
JER|48|12|看哪，日子将到，我必差倒酒的到它那里去，将它倒出来；他们要倒空器皿，打碎坛子。这是耶和华说的。
JER|48|13|摩押 必因 基抹 羞愧，像 以色列 家因倚靠 伯特利 羞愧一样。
JER|48|14|你们怎么说： “我们是勇士，是会打仗的壮士”呢？
JER|48|15|摩押 变为废墟， 敌人上去占它的城镇。 它精良的壮丁都下去遭杀戮； 这是名为万军之耶和华的君王说的。
JER|48|16|摩押 的灾殃临近， 灾难速速来到。
JER|48|17|凡在它四围的和认识它名的， 都要为它悲伤，说： 那结实的杖和美好的棍， 竟然折断了！
JER|48|18|底本 的居民哪， 要从你荣耀的座位上下来， 坐着忍受干渴； 因毁灭 摩押 的人上来攻击你， 毁坏了你的堡垒。
JER|48|19|住 亚罗珥 的啊， 要站在道路的边上观望， 问逃跑的男人和逃脱的女人说： “发生了什么事呢”？
JER|48|20|摩押 因毁坏蒙羞； 你们要哀号呼喊， 要在 亚嫩 报告： “ 摩押 已成废墟！”
JER|48|21|审判临到平原之地的 何伦 、 雅杂 、 米法押 、
JER|48|22|底本 、 尼波 、 伯．低比拉太音 、
JER|48|23|基列亭 、 伯．迦末 、 伯．米恩 、
JER|48|24|加略 、 波斯拉 和 摩押 地远近所有的城镇。
JER|48|25|摩押 的角砍断了，膀臂折断了。这是耶和华说的。
JER|48|26|你们要使 摩押 沉醉，因它向耶和华夸大。它要在自己所吐之物中打滚，又要被人嗤笑。
JER|48|27|以色列 不是你的笑柄吗？它难道是在贼中被逮到，使你每逢提到它就摇头的吗？
JER|48|28|摩押 的居民哪， 要离开城镇，住在山崖里， 像鸽子在峡谷口上搭窝。
JER|48|29|我们听闻 摩押 人的骄傲， 极其骄傲； 他们自高、自傲、 自我狂妄、居心自大。
JER|48|30|我知道他们的愤怒是虚空的， 他们夸大的话一无所成。 这是耶和华说的。
JER|48|31|因此，我要为 摩押 哀号， 为 摩押 全地呼喊； 人必为 吉珥．哈列设 人叹息。
JER|48|32|西比玛 的葡萄树啊，我为你哀哭， 甚于 雅谢 人的哀哭。 你的枝子蔓延过海， 直伸到 雅谢海 。 那行毁灭的已经临到你夏天的果子和葡萄。
JER|48|33|肥田和 摩押 地的欢喜快乐都被夺去， 我使酒池不再流出酒来， 无人踹酒欢呼； 呼喊的声音不再是欢呼。
JER|48|34|有哀声从 希实本 达到 以利亚利 ，他们发的哀声达到 雅杂 ；从 琐珥 达到 何罗念 ，达到 伊基拉．施利施亚 ，因为 宁林 的水必然干涸。
JER|48|35|我必在 摩押 地使那在丘坛献祭的，和那向他的神明烧香的都灭绝了。这是耶和华说的。
JER|48|36|因此，我的心为 摩押 哀鸣如箫，我的心为 吉珥．哈列设 人哀哭； 摩押 人所得的财物都毁灭了。
JER|48|37|各人头上光秃，胡须剪短，手有划伤，腰束麻布。
JER|48|38|在 摩押 的各房顶上和街市上到处有人哀哭，因我打碎 摩押 ，好像打碎无人喜爱的器皿。这是耶和华说的。
JER|48|39|打得粉碎了！他们要哀号了！ 摩押 要羞愧转背了！这样， 摩押 必受四围的人嗤笑惊骇。
JER|48|40|耶和华如此说： 看哪，仇敌必如鹰展翅快飞， 攻击 摩押 。
JER|48|41|加略 被攻取，堡垒也被占据。 到那日， 摩押 的勇士心中疼痛如临产的妇人。
JER|48|42|摩押 必被毁灭，不再成国， 因它向耶和华夸大。
JER|48|43|摩押 的居民哪， 惊吓、陷阱、罗网都临近你。 这是耶和华说的。
JER|48|44|躲过惊吓的必坠入陷阱， 逃离陷阱的又被罗网缠住， 因我必使惩罚之年临到 摩押 。 这是耶和华说的。
JER|48|45|逃难的人站在 希实本 的荫下，筋疲力尽， 因为有火从 希实本 发出， 有火焰出自 西宏 ， 烧尽 摩押 的鬓角和闹哄人的头顶。
JER|48|46|摩押 啊，你有祸了！ 属 基抹 的百姓灭亡了！ 因你的儿子都被掳去， 你的女儿也被掳去。
JER|48|47|到末后，我却要使 摩押 被掳的人归回。 摩押 受审判的话到此为止。 这是耶和华说的。
JER|49|1|论 亚扪 人。 耶和华如此说： 以色列 没有儿子吗？ 没有后嗣吗？ 米勒公 为何承受 迦得 为业呢？ 属它的百姓为何住其中的城镇呢？
JER|49|2|看哪，日子将到，我必使人听见打仗的喊声， 攻击 亚扪 人所住的 拉巴 的喊声。 拉巴 要成为废墟， 属它的乡镇 要被火焚烧。 这是耶和华说的。 先前承受 以色列 为业的， 此时 以色列 倒要承受他们为业。 这是耶和华说的。
JER|49|3|希实本 哪，要哀号， 因为 爱 地已成荒地。 拉巴 的乡镇哪，要呼喊， 以麻布束腰； 要哭号，在篱笆中往来奔跑； 因 米勒公 和它的祭司、 官长要一同被掳去。
JER|49|4|背道的民 哪， 你为何因有山谷， 因有水流的山谷夸耀呢？ 为何倚靠自己的财宝，说： “谁能来到我们这里呢？”
JER|49|5|万军之主耶和华说： 看哪，我要使惊吓从四围的邻邦临到你们； 你们必被赶出， 各人一直往前， 无人收容难民。
JER|49|6|但后来，我却要使被掳的 亚扪 人归回。这是耶和华说的。
JER|49|7|论 以东 。 万军之耶和华如此说： 提幔 不再有智慧了吗？ 聪明人的谋略都用尽了吗？ 他们的智慧尽归无有了吗？
JER|49|8|底但 的居民哪，要转身逃跑， 住在深密处； 因为我惩罚 以扫 的时候， 必使灾殃临到他。
JER|49|9|摘葡萄的若来到你那里， 岂不留下几串吗？ 贼若夜间来到， 岂不是只毁坏他们要毁坏的吗？
JER|49|10|我却使 以扫 赤裸， 暴露他的藏身处； 他不能隐藏自己。 他的后裔、弟兄、邻舍全都灭绝， 他也归于无有。
JER|49|11|你撇下孤儿，我必保全他们的性命； 你的寡妇可以倚靠我。
JER|49|12|耶和华如此说：“看哪，既然原不该喝那杯的一定要喝，你能免去惩罚吗？必不能免，一定要喝！
JER|49|13|我指着自己起誓， 波斯拉 必令人惊骇、受羞辱、被诅咒，并且全然荒废。它所有的城镇都要永远成为废墟。这是耶和华说的。”
JER|49|14|我从耶和华那里听见消息， 有使者被差往列国去，说： “你们要聚集前来攻击 以东 ， 要起来争战。”
JER|49|15|看哪，我使你在列国中为最小， 在世人中被藐视。
JER|49|16|住在山穴中盘据山顶的啊， 你被自己的声势与心中的狂傲所蒙蔽； 你虽如大鹰高高搭窝， 我却要从那里拉你下来。 这是耶和华说的。
JER|49|17|以东 必令人惊骇；凡经过的人都惊骇，又因它一切的灾祸嗤笑。
JER|49|18|耶和华说：它要像 所多玛 、 蛾摩拉 和邻近的城镇一样倾覆，必无人住在那里，也无人在其中寄居。
JER|49|19|看哪，就像狮子从 约旦河 边的丛林上来，攻击坚固的居所，我要在转眼之间使 以东 人逃跑，离开这地。我拣选谁，就派谁治理这地。谁能像我呢？谁能召我出庭呢？ 有哪一个牧人能在我面前站得住呢？
JER|49|20|你们要听耶和华攻击 以东 所定的计划和他攻击 提幔 居民所定的旨意。他们羊群当中微弱的定要被拖走，他们的草场定要变为荒凉。
JER|49|21|因他们仆倒的声音，地就震动，哀号的声音传到 红海 那里。
JER|49|22|看哪，仇敌必如大鹰飞起，展开翅膀攻击 波斯拉 。到那日， 以东 的勇士心中疼痛如临产的妇人。
JER|49|23|论 大马士革 。 哈马 和 亚珥拔 蒙羞， 因为他们听见凶恶的消息就融化； 焦虑像海浪汹涌，不得平静。
JER|49|24|大马士革 发软，转身逃跑； 战兢将它捉住， 痛苦忧愁将它抓住， 如临产的妇人一样。
JER|49|25|我所喜乐受称赞的城， 怎能被撇弃 呢？
JER|49|26|它的壮丁必仆倒在街上， 当那日，战士全都静默无声。 这是万军之耶和华说的。
JER|49|27|我必用火点燃 大马士革 的城墙， 烧灭 便．哈达 的宫殿。
JER|49|28|论 巴比伦 王 尼布甲尼撒 所攻打的 基达 和 夏琐 诸国。 耶和华如此说： 迦勒底 人哪，起来上 基达 去， 毁灭东方人。
JER|49|29|人要夺去他们的帐棚和羊群， 人要带走他们的幔子、一切器皿，和骆驼，占为己有。 人向他们喊着说： 四围都有惊吓。
JER|49|30|夏琐 的居民哪，要逃奔远方， 住在深远之处； 因为 巴比伦 王 尼布甲尼撒 设计谋害你们， 起意攻击你们。 这是耶和华说的。
JER|49|31|迦勒底 人哪，起来！ 上到安逸无虑的国民那里去， 他们是无门无闩、单独居住的。 这是耶和华说的。
JER|49|32|他们的骆驼必成为掠物， 他们众多的牲畜必成为掳物。 我要将剃鬓发的人分散四方 ， 使灾殃从四围临到他们。 这是耶和华说的。
JER|49|33|夏琐 必成为野狗的住处， 永远荒废； 无人住在那里， 也无人在其中寄居。
JER|49|34|犹大 王 西底家 登基的时候，耶和华论 以拦 的话临到 耶利米 先知，说：
JER|49|35|“万军之耶和华如此说：看哪，我必折断 以拦 人的弓，那是他们战斗的主力。
JER|49|36|我要使风从天的四方刮来，临到 以拦 ，将他们分散四方。 以拦 被赶散的人没有一国不到的。
JER|49|37|我必使 以拦 人在仇敌和寻索其命的人面前惊惶；我也必使灾祸，就是我的烈怒临到他们，又必使刀剑追杀他们，直到将他们灭尽。这是耶和华说的。
JER|49|38|我要在 以拦 设立我的宝座，在那里除灭君王和官长。这是耶和华说的。
JER|49|39|“到末后，我却要使被掳的 以拦 人归回。这是耶和华说的。”
JER|50|1|以下是耶和华藉 耶利米 先知论 巴比伦 和 迦勒底 人之地所说的话。
JER|50|2|你们要在万国中传扬，宣告， 竖立大旗； 要宣告，不可隐瞒，说： “ 巴比伦 被攻取， 彼勒 蒙羞， 米罗达 惊惶。 巴比伦 的神像都蒙羞， 它的偶像都惊惶。”
JER|50|3|因有一国从北方上来攻击它，使它的地荒凉，无人居住，连人带牲畜都逃走了。
JER|50|4|在那日、在那时， 以色列 人要和 犹大 人同来，随走随哭，寻求耶和华－他们的上帝。这是耶和华说的。
JER|50|5|他们要问到 锡安 之路，又面向那里，说：“来吧，他们要 在永不被遗忘的约中与耶和华联合。”
JER|50|6|我的百姓成了失丧的羊，牧人使他们走迷了路，转入丛山之间。他们从大山走到小山，竟忘了自己安歇之处。
JER|50|7|凡遇见他们的，就把他们吞灭。敌人说：“我们不算有罪；因他们得罪了那可作真正 居所的耶和华，就是他们祖先所仰望的耶和华。”
JER|50|8|“你们要逃离 巴比伦 ，要离开 迦勒底 人之地，像走在羊群前面的公山羊。
JER|50|9|看哪，因我必激起大国联盟，带领他们从北方来攻击 巴比伦 ，他们要摆阵攻击它，它必在那里被攻取。他们的箭好像善射 勇士的箭，绝不徒然返回。
JER|50|10|迦勒底 要成为掠物，凡掳掠它的都必心满意足。这是耶和华说的。”
JER|50|11|抢夺我产业的啊， 你们因欢喜快乐， 像踹谷 嬉戏的母牛犊， 又像发嘶声的壮马。
JER|50|12|你们的母亲极其抱愧， 生你们的必然蒙羞。 看哪，她要列在诸国之末， 成为旷野、旱地、沙漠；
JER|50|13|因耶和华的愤怒， 巴比伦 必无人居住， 全然荒凉， 凡经过的都要受惊骇， 又因它所遭的灾殃嗤笑。
JER|50|14|所有拉弓的啊，要在 巴比伦 的四围摆阵， 射箭攻击它， 不用爱惜箭枝， 因为它得罪了耶和华。
JER|50|15|要在它四围呐喊： “它已经投降， 堡垒坍塌了， 城墙拆毁了！” 这是耶和华所报的仇。 你们要向它报仇； 它怎样待人，你们也要怎样待它。
JER|50|16|你们要将 巴比伦 撒种的 和收割时拿镰刀的全都剪除。 他们各人因躲避欺压的刀剑， 必归回本族，逃到本土。
JER|50|17|以色列 是打散的羊，被狮子赶散。首先是 亚述 王将他吞灭，末后是 巴比伦 王 尼布甲尼撒 折断他的骨头。
JER|50|18|所以万军之耶和华－ 以色列 的上帝如此说：“看哪，我必惩罚 巴比伦 王和他的地，像我从前惩罚 亚述 王一样。
JER|50|19|我必领 以色列 回他自己的草场，他要在 迦密 和 巴珊 吃草，又在 以法莲 山上和 基列 境内得以饱足。
JER|50|20|在那日、在那时，你寻找 以色列 的罪孽，一无所有；寻找 犹大 的罪恶，也无所得；因为我所留下的人，我必赦免。这是耶和华说的。”
JER|50|21|你要上去攻击 米拉大翁 之地， 又攻击 比割 的居民。 将他们追杀灭尽， 照我所吩咐你的一切去做。 这是耶和华说的。
JER|50|22|境内有打仗和大毁灭的响声。
JER|50|23|全地的大锤竟然砍断破坏！ 巴比伦 在列国中竟然荒凉！
JER|50|24|巴比伦 哪，我为你设下罗网， 你被缠住，竟不自觉。 你被寻着，也被捉住， 因为你对抗耶和华。
JER|50|25|耶和华已经打开军械库， 拿出他恼恨的兵器； 这是万军之主耶和华 在 迦勒底 人之地要做的事。
JER|50|26|你们要从极远的边界前来攻击它 ， 要开它的仓廪， 将它堆起如高堆， 毁灭净尽，丝毫不留。
JER|50|27|要杀它一切的牛犊， 使它们下去遭杀戮。 他们有祸了， 因为他们的日子，就是他们受罚的时刻已经来到。
JER|50|28|从 巴比伦 之地逃出来的难民，在 锡安 扬声宣告耶和华－我们的上帝要报仇，为他的圣殿报仇。
JER|50|29|你们要招集一切弓箭手来攻击 巴比伦 ，在 巴比伦 四围安营，不容一人逃脱。要照着它所做的报应它；它怎样待人，你们也要怎样待它，因为它向耶和华－ 以色列 的圣者狂傲。
JER|50|30|所以它的壮丁必仆倒在街上。当那日，它的士兵全都静默无声。这是耶和华说的。
JER|50|31|“看哪，你这狂傲的啊，我与你为敌， 因为你的日子， 我惩罚你的时刻已经来到。 这是万军之主耶和华说的。
JER|50|32|狂傲的必绊跌仆倒，无人扶起。 我必用火点燃他的城镇， 将他四围所有的尽行烧灭。”
JER|50|33|万军之耶和华如此说：“ 以色列 人和 犹大 人一同受欺压；凡掳掠他们的都紧紧抓住他们，不肯释放。
JER|50|34|他们的救赎主大有能力，万军之耶和华是他的名。他必定为他们伸冤，使全地得享平静；他却要搅扰 巴比伦 的居民。”
JER|50|35|有刀剑临到 迦勒底 人和 巴比伦 的居民， 临到它的领袖与智慧人。 这是耶和华说的。
JER|50|36|有刀剑临到矜夸的人， 他们就变为愚昧； 有刀剑临到它的勇士， 他们就惊惶。
JER|50|37|有刀剑临到它的马匹、战车， 和其中混居的各族， 他们变成与妇女一样； 有刀剑临到它的宝物， 宝物就被抢夺。
JER|50|38|有干旱 临到它的众水， 它们就必干涸； 因为这是雕刻偶像之地， 人因偶像颠狂 。
JER|50|39|所以野兽和土狼必住在那里，鸵鸟也住在其中，永远无人居住，世世代代无人定居。
JER|50|40|巴比伦 要像上帝所倾覆的 所多玛 、 蛾摩拉 和邻近的城镇一样，必无人住在那里，也无人在其中寄居。这是耶和华说的。
JER|50|41|看哪，有一民族从北方而来， 有一大国和许多君王被激起，从地极来到。
JER|50|42|他们拿弓和枪， 性情残忍，毫不留情； 他们的声音像海浪澎湃。 巴比伦 啊， 他们骑着马， 如上战场的人摆列队伍， 要攻击你。
JER|50|43|巴比伦 王听见他们的风声， 手就发软， 痛苦将他抓住， 仿佛临产的妇人疼痛一般。
JER|50|44|“看哪，就像狮子从 约旦河 边的丛林上来，攻击坚固的居所，我要在转眼之间使 迦勒底 人逃跑，离开这地。我拣选谁，就派谁治理这地。谁能像我呢？谁能召我出庭呢？有哪一个牧人能在我面前站得住呢？
JER|50|45|你们要听耶和华攻击 巴比伦 所定的计划和他攻击 迦勒底 人之地所定的旨意。他们羊群当中微弱的定要被拖走，他们的草场定要变为荒凉。
JER|50|46|因 巴比伦 被攻下的声音，地就震动，人在列国都听见呼喊的声音。”
JER|51|1|耶和华如此说： 看哪，我必刮起毁灭的风， 攻击 巴比伦 和住在 立加米 的人。
JER|51|2|我要差陌生人 来到 巴比伦 ， 他们要簸扬它，使它的地空无一物。 在它遭祸的日子， 他们要四围攻击它。
JER|51|3|不要叫拉弓的拉弓， 不要叫他佩戴盔甲 ； 不要怜惜 巴比伦 的壮丁， 要灭尽它的全军。
JER|51|4|他们必在 迦勒底 人之地被杀仆倒， 在 巴比伦 的街市上被刺透。
JER|51|5|以色列 和 犹大 境内虽然充满违背 以色列 圣者的罪， 却没有被他的上帝－万军之耶和华所遗弃。
JER|51|6|你们要奔逃，离开 巴比伦 ， 各救自己的性命！ 不要陷在它的罪孽中一同灭亡， 因为这是耶和华报仇的时刻， 他必向 巴比伦 施行报应。
JER|51|7|巴比伦 素来是耶和华手中的金杯， 使全地沉醉， 列国喝了它的酒就颠狂。
JER|51|8|巴比伦 忽然倾覆毁坏； 要为它哀号， 拿乳香来止它的疼痛， 或者可以治好。
JER|51|9|我们想医治 巴比伦 ， 它却未获痊愈。 离开它吧！让我们各人归回本国， 因为它受的审判通于上天，达到穹苍。
JER|51|10|耶和华已经彰显出我们的义。 来吧！我们要在 锡安 传扬耶和华－我们上帝的作为。
JER|51|11|你们要磨尖箭头， 抓住盾牌。 论到 巴比伦 ，耶和华定意要毁灭它，所以激起 玛代 君王的心；这是耶和华报仇，为他的圣殿报仇。
JER|51|12|你们要竖立大旗， 攻击 巴比伦 的城墙； 要坚固了望台， 派定守望的设下埋伏； 因为耶和华指着 巴比伦 居民所说的， 他不但这样定意，也已成就。
JER|51|13|住在众水之上多有财宝的啊， 你的结局已到！ 你贪婪之量已满盈 ！
JER|51|14|万军之耶和华指着自己起誓说： 我必使人遍满各处像蝗虫一样， 他们必呐喊攻击你。
JER|51|15|耶和华以能力创造大地， 以智慧建立世界， 以聪明铺张穹苍。
JER|51|16|他一出声，天上就有众水澎湃； 他使云雾从地极上腾， 造电随雨而闪， 从仓库中吹出风来。
JER|51|17|人人都如同畜牲，毫无知识； 银匠都因偶像羞愧， 他所铸的偶像本为虚假， 它们里面并无气息。
JER|51|18|它们都是虚无的， 是迷惑人的东西， 到它们受罚的时刻必被除灭。
JER|51|19|雅各 所得的福分不是这样， 因主 是那创造万有的， 以色列 是他产业的支派， 万军之耶和华是他的名。
JER|51|20|你是我争战的斧子和打仗的兵器。 我要用你打碎列邦， 毁灭列国；
JER|51|21|用你打碎马和骑马的， 打碎战车和坐在其上的；
JER|51|22|用你打碎男人和女人， 打碎老人和少年， 打碎壮丁和少女；
JER|51|23|用你打碎牧人和他的羊群， 打碎农夫和他的一对耕牛， 打碎省长和官员。
JER|51|24|我必在你们眼前报复 巴比伦 人和 迦勒底 居民在 锡安 所做的一切恶事。这是耶和华说的。
JER|51|25|行毁灭的山，看哪，我与你为敌， 你毁灭全地， 我必伸手攻击你， 将你从山岩滚下去， 使你成为烧毁了的山。 这是耶和华说的。
JER|51|26|人必不从你那里取石头为房角石， 也不取石头来作根基， 因为你必永远荒废。 这是耶和华说的。
JER|51|27|你们要在境内竖立大旗， 在列邦中吹角， 使列邦预备攻击 巴比伦 。 要招集 亚拉腊 、 米尼 、 亚实基拿 各国前来攻击它， 派将军攻击它， 使马匹上来如粗暴的蝗虫；
JER|51|28|使列邦和 玛代 君王，省长和官员， 他们所管的全地，都预备攻击它。
JER|51|29|地必震动而移转； 因耶和华向 巴比伦 旨意已确定， 要使 巴比伦 土地荒凉，无人居住。
JER|51|30|巴比伦 的勇士停止争战， 躲在堡垒之中。 他们的力气耗尽， 他们变成与妇女一样。 巴比伦 的住处焚烧， 门闩都折断了。
JER|51|31|通报的彼此相遇， 送信的彼此相遇， 报告 巴比伦 王， 城的四方都被攻下了，
JER|51|32|渡口被占据了， 芦苇被火焚烧， 战士都惊慌。
JER|51|33|万军之耶和华－ 以色列 的上帝如此说： 巴比伦 好像踹谷的禾场； 再过片时，它收割的时候就到了。
JER|51|34|巴比伦 王 尼布甲尼撒 吞灭我，压碎我， 使我成为空器皿。 他如大鱼将我吞下， 以我的美物充满他的肚腹， 又把我赶出去。
JER|51|35|锡安 的居民要说： 愿我和我骨肉之亲所受的残暴 归给 巴比伦 。 耶路撒冷 人要说： 愿我们所流的血 归给 迦勒底 的居民。
JER|51|36|所以，耶和华如此说： 看哪，我必为你伸冤，为你报仇； 我必使 巴比伦 的海枯竭， 使它的泉源干涸。
JER|51|37|巴比伦 必成为废墟， 为野狗的住处， 令人惊骇、嗤笑， 并且无人居住。
JER|51|38|他们要像少壮狮子一同咆哮， 像小狮子吼叫。
JER|51|39|他们食欲一来的时候， 我必为他们摆设酒席， 使他们沉醉，好叫他们快乐； 他们睡了长觉，永不醒起。 这是耶和华说的。
JER|51|40|我必使他们像羔羊、 像公绵羊和公山羊被牵去宰杀。
JER|51|41|示沙克 竟然被攻取！ 全地所称赞的被占据！ 巴比伦 在列国中竟然变为荒凉！
JER|51|42|海水涨起，漫过 巴比伦 ； 澎湃的海浪遮盖了它。
JER|51|43|它的城镇变废墟， 地变干旱，成为沙漠， 成为无人居住、 无人经过之地。
JER|51|44|我要惩罚 巴比伦 的 彼勒 ， 使它吐出所吞之物。 列国必不再流归到它那里， 巴比伦 的城墙也必坍塌。
JER|51|45|我的子民哪，你们要离开 巴比伦 ！ 各人逃命，躲避耶和华的烈怒。
JER|51|46|不要因境内所听见的风声 心惊胆怯或惧怕； 因为这年有风声传来， 那年也有风声传来； 境内有残暴的事， 官长攻击官长。
JER|51|47|所以，看哪，日子将到， 我必惩罚 巴比伦 雕刻的偶像。 它的全地必然抱愧， 它被杀的人必仆倒在其上。
JER|51|48|那时，天地和其中所有的， 必因 巴比伦 欢呼， 因为行毁灭的要从北方来到它那里。 这是耶和华说的。
JER|51|49|巴比伦 要因 以色列 被杀的人而仆倒， 正如全地被刺杀的人是因 巴比伦 仆倒一般。
JER|51|50|你们躲避刀剑的要快走， 不要站住！ 要在远方怀念耶和华， 心中追想 耶路撒冷 。
JER|51|51|我们听见辱骂就蒙羞，满面惭愧， 因为外邦人进入耶和华殿的圣所。
JER|51|52|所以，看哪，日子将到， 我必惩罚 巴比伦 雕刻的偶像， 在全境内到处都有刺伤的人在呻吟。 这是耶和华说的。
JER|51|53|巴比伦 虽升到天上， 虽使它坚固的高处更坚固， 我也要差毁灭者到它那里。 这是耶和华说的。
JER|51|54|有哀号的声音从 巴比伦 出来， 有大毁灭从 迦勒底 人之地而来。
JER|51|55|耶和华使 巴比伦 变为废墟， 使其中喧哗的大声灭绝。 仇敌仿佛众水， 波浪澎湃，发出响声；
JER|51|56|这是行毁灭的临到 巴比伦 。 巴比伦 的勇士被捉住， 他们的弓折断了； 因为耶和华是施行报应的上帝， 他必施行报应。
JER|51|57|我必使 巴比伦 的领袖、 智慧人、省长、官员和勇士都喝醉， 使他们永远沉睡，不再醒起。 这是名为万军之耶和华的君王说的。
JER|51|58|万军之耶和华如此说： 巴比伦 宽阔的城墙要夷为平地， 它高大的城门必被火焚烧。 万民所劳碌的必致虚空， 万族所劳碌的被火焚烧， 他们都必困乏。
JER|51|59|犹大 王 西底家 在位第四年， 玛西雅 的孙子， 尼利亚 的儿子 西莱雅 与王同去 巴比伦 ， 西莱雅 是王宫的大臣， 耶利米 先知有话吩咐他。
JER|51|60|耶利米 把一切要临到 巴比伦 的灾祸，就是论到 巴比伦 的这一切话，写在一书卷上。
JER|51|61|耶利米 对 西莱雅 说：“你到了 巴比伦 ，务要宣读这一切话，
JER|51|62|说：‘耶和华啊，你曾论到这地方说：要剪除它，不再有人与牲畜居住此地，必永远荒凉。’
JER|51|63|你读完这书卷，就要把一块石头拴在其上，投入 幼发拉底河 中，
JER|51|64|说：‘ 巴比伦 因耶和华所要降与它的灾祸，必如此沉下去，不再浮起来，百姓也必困乏。’” 耶利米 的话到此为止。
JER|52|1|西底家 登基的时候年二十一岁，在 耶路撒冷 作王十一年。他母亲名叫 哈慕她 ，是 立拿 人 耶利米 的女儿。
JER|52|2|西底家 行耶和华眼中看为恶的事，像 约雅敬 所做的一切。
JER|52|3|因此，耶和华向 耶路撒冷 和 犹大 发怒，以致把他们从自己面前赶出去。 西底家 背叛 巴比伦 王，
JER|52|4|他作王第九年十月初十， 巴比伦 王 尼布甲尼撒 率领全军前来攻击 耶路撒冷 ，对着城安营，四围筑堡垒攻城，
JER|52|5|城被围困，直到 西底家 王十一年。
JER|52|6|四月初九，城里的饥荒非常严重，当地的百姓都没有粮食。
JER|52|7|城被攻破，士兵全都在夜间从靠近王园两城墙中间的门逃跑出城； 迦勒底 人正在四围攻城，他们就往 亚拉巴 逃去。
JER|52|8|迦勒底 的军队追赶 西底家 王，在 耶利哥 的平原追上他。他的全军都离开他溃散了。
JER|52|9|迦勒底 人就拿住王，带他到 哈马 地 利比拉 的 巴比伦 王那里； 巴比伦 王就判他的罪。
JER|52|10|巴比伦 王在 西底家 眼前杀了他的儿女，又在 利比拉 杀了 犹大 全体的官长，
JER|52|11|并且挖了 西底家 的眼睛，用铜链锁着他，带到 巴比伦 去，将他囚在监里，直到他死的日子。
JER|52|12|巴比伦 王 尼布甲尼撒 十九年五月初十，在 巴比伦 王面前侍立的 尼布撒拉旦 护卫长进入 耶路撒冷 ，
JER|52|13|他焚烧了耶和华的殿、王宫和 耶路撒冷 的房屋；用火焚烧所有大户人家的房屋。
JER|52|14|跟随护卫长的 迦勒底 全军拆毁了 耶路撒冷 四围的城墙。
JER|52|15|那时 尼布撒拉旦 护卫长将百姓中最穷的和城里所剩下的百姓，并那些投降 巴比伦 王的人，以及剩下的工匠，都掳去了。
JER|52|16|但 尼布撒拉旦 护卫长留下一些当地最穷的人，叫他们修整葡萄园，耕种田地。
JER|52|17|耶和华殿的铜柱并殿内的盆座和铜海， 迦勒底 人都打碎了，把那些铜运到 巴比伦 去；
JER|52|18|他们又带走锅、铲子、钳子、盘子、勺子，和供奉用的一切铜器；
JER|52|19|杯、火盆、碗、锅、灯台、勺子、酒杯，无论金的银的，护卫长都带走了；
JER|52|20|还有 所罗门 为耶和华殿所造的两根柱子、一面铜海，并座下的十二只铜牛，这些器皿的铜多得无法可秤。
JER|52|21|至于柱子，这一根柱子高十八肘，厚四指，周围十二肘，中间是空的；
JER|52|22|柱上有铜顶，每个铜顶高五肘；铜顶的周围有网子和石榴，也都是铜的。另一根柱子与此相同，也有石榴。
JER|52|23|柱子四面有九十六个石榴，在网子周围，总共有一百个石榴。
JER|52|24|护卫长拿住 西莱雅 大祭司、 西番亚 副祭司和门口的三个守卫，
JER|52|25|又从城中拿住一个管理士兵的官 ，并在城里找到王面前的七个亲信，和召募当地百姓之将军的书记官，以及在城中找到的六十个当地百姓。
JER|52|26|尼布撒拉旦 护卫长把这些人带到 利比拉 的 巴比伦 王那里。
JER|52|27|巴比伦 王击杀他们，在 哈马 地的 利比拉 把他们处死。这样， 犹大 人就被掳去离开本地。
JER|52|28|这是 尼布甲尼撒 所掳百姓的数目：他在位第七年掳去 犹大 人三千零二十三人；
JER|52|29|尼布甲尼撒 十八年从 耶路撒冷 掳去八百三十二人；
JER|52|30|尼布甲尼撒 二十三年， 尼布撒拉旦 护卫长掳去 犹大 人七百四十五人；共有四千六百人。
JER|52|31|巴比伦 王 以未．米罗达 作王的元年，就是 犹大 王 约雅斤 被掳后三十七年十二月二十五日，他使 犹大 王 约雅斤 抬起头来，提他出监，
JER|52|32|对他说好话，使他的位高过与他一同被掳、在 巴比伦 众王的位；
JER|52|33|又给他脱了囚服，使他终身常在 巴比伦 王面前吃饭。
JER|52|34|巴比伦 王赐给他日常需用的食物，日日一份，终身都是这样，直到他死的日子。
