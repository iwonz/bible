GEN|1|1|起初，上帝創造天地。
GEN|1|2|地是空虛混沌，深淵上面一片黑暗；上帝的靈 運行在水面上。
GEN|1|3|上帝說：「要有光」，就有了光。
GEN|1|4|上帝看光是好的，於是上帝就把光和暗分開。
GEN|1|5|上帝稱光為「晝」，稱暗為「夜」。有晚上，有早晨，這是第一日。
GEN|1|6|上帝說：「眾水之間要有穹蒼，把水和水分開。」
GEN|1|7|上帝就造了穹蒼，把穹蒼以下的水和穹蒼以上的水分開。事就這樣成了。
GEN|1|8|上帝稱穹蒼為「天」。有晚上，有早晨，這是第二日。
GEN|1|9|上帝說：「天下面的水要聚集在一處，使乾地露出來。」事就這樣成了。
GEN|1|10|上帝稱乾地為「地」，稱聚集在一起的水為「海」。上帝看為好的。
GEN|1|11|上帝說：「地要長出植物，就是含種子的五穀菜蔬，和會結果子、果子裏有種子的樹，在地上各從其類。」事就這樣成了。
GEN|1|12|於是地長出了植物：含種子的五穀菜蔬，各從其類；會結果子、果子裏有種子的樹，各從其類。上帝看為好的。
GEN|1|13|有晚上，有早晨，這是第三日。
GEN|1|14|上帝說：「天上要有光體來分晝夜，讓它們作記號，定季節、日子、年份，
GEN|1|15|它們要在天空發光，照在地上。」事就這樣成了。
GEN|1|16|於是上帝造了兩個大光體，大的管晝，小的管夜，又造了星辰。
GEN|1|17|上帝把這些光體擺列在天空，照在地上，
GEN|1|18|管理晝夜，分別光暗。上帝看為好的。
GEN|1|19|有晚上，有早晨，這是第四日。
GEN|1|20|上帝說：「水要滋生眾多有生命之物；要有鳥飛在地面以上，天空之中。」
GEN|1|21|上帝就創造了大魚和在水裏滋生的各樣活動的生物，各從其類，以及各樣有翅膀的鳥，各從其類。上帝看為好的。
GEN|1|22|上帝就賜福給這一切，說：「要繁殖增多，充滿在海的水裏；飛鳥也要在地上增多。」
GEN|1|23|有晚上，有早晨，這是第五日。
GEN|1|24|上帝說：「地要生出有生命之物，各從其類，就是牲畜、爬行動物、地上的走獸，各從其類。」事就這樣成了。
GEN|1|25|於是上帝造了地上的走獸，各從其類；牲畜，各從其類；和地上一切的爬行動物，各從其類。上帝看為好的。
GEN|1|26|上帝說：「我們要照著我們的形像，按著我們的樣式造人，使他們管理海裏的魚、天空的鳥、地上的牲畜和全地，以及地上爬的一切爬行動物。」
GEN|1|27|上帝就照著他的形像創造人，照著上帝的形像創造他們 ；他創造了他們，有男有女。
GEN|1|28|上帝賜福給他們，上帝對他們說：「要生養眾多，遍滿這地，治理它；要管理海裏的魚、天空的鳥和地上各樣活動的生物。」
GEN|1|29|上帝說：「看哪，我把全地一切含種子的五穀菜蔬和一切會結果子、果子裏有種子的樹，都賜給你們；這些都可作食物。
GEN|1|30|至於地上一切的走獸、天空一切的飛鳥，並一切在地上爬行的，有生命的動物，我把綠色植物賜給牠們作食物。」事就這樣成了。
GEN|1|31|上帝看一切所造的，看哪，都非常好。有晚上，有早晨，這是第六日。
GEN|2|1|天和地，以及萬象都完成了。
GEN|2|2|到第七日，上帝已經完成了造物之工，就在第七日安息了，歇了他所做一切的工。
GEN|2|3|上帝賜福給第七日，將它分別為聖，因為在這日，上帝安息了，歇了他所做一切創造的工。
GEN|2|4|這就是天地創造的來歷。 在耶和華上帝造地和天的時候，
GEN|2|5|地上還沒有田野的草木，田間的菜蔬還沒有長出來，因為耶和華上帝還沒有降雨在地上，也沒有人耕種土地。
GEN|2|6|但是，有霧氣從地上騰，滋潤整個土地的表面。
GEN|2|7|耶和華上帝用地上的塵土造人，將生命之氣吹進他的鼻孔，這人就成了有靈的活人 。
GEN|2|8|耶和華上帝在東方的 伊甸 栽了一個園子，把所造的人安置在那裏。
GEN|2|9|耶和華上帝使各樣的樹從土地裏長出來，可以悅人的眼目，好作食物。園子當中有生命樹和知善惡的樹 。
GEN|2|10|有一條河從 伊甸 流出來，滋潤那園子，從那裏分成四個源頭：
GEN|2|11|第一條名叫 比遜 ，它環繞 哈腓拉 全地，在那裏有金子。
GEN|2|12|那地的金子很好，在那裏也有珍珠 和紅瑪瑙。
GEN|2|13|第二條河名叫 基訓 ，它環繞 古實 全地。
GEN|2|14|第三條河名叫 底格里斯 ，它流到 亞述 的東邊。第四條河就是 幼發拉底 。
GEN|2|15|耶和華上帝把那人安置在 伊甸園 ，讓他耕耘看管。
GEN|2|16|耶和華上帝吩咐那人說：「園中各樣樹上所出的，你可以隨意吃，
GEN|2|17|只是知善惡的樹所出的，你不可吃，因為你吃它的日子必定死！」
GEN|2|18|耶和華上帝說：「那人單獨一個不好，我要為他造一個配偶幫助他。」
GEN|2|19|耶和華上帝用泥土造了野地各樣的走獸和天空各樣的飛鳥，都帶到那人面前，看他叫甚麼。那人怎樣叫各樣的動物，那就是牠的名字。
GEN|2|20|那人就給一切牲畜、天空的飛鳥和野地各樣的走獸都起了名。只是 亞當 沒有找到配偶幫助他。
GEN|2|21|耶和華上帝使他沉睡，他就睡了；於是取下他的一根肋骨，又在原處把肉合起來。
GEN|2|22|耶和華上帝就用那人身上所取的肋骨造了一個女人，帶她到那人面前。
GEN|2|23|那人說： 「這正是我骨中的骨， 肉中的肉， 可以稱她為女人， 因為她是從男人身上取出來的。」
GEN|2|24|因此，人要離開父母，與妻子結合，二人成為一體。
GEN|2|25|當時夫妻二人赤身露體，並不覺得羞恥。
GEN|3|1|耶和華上帝所造的，惟有蛇比田野一切的走獸更狡猾。蛇對女人說：「上帝豈是真說，你們不可吃園中任何樹上所出的嗎？」
GEN|3|2|女人對蛇說：「園中樹上的果子，我們都可以吃；
GEN|3|3|只是園子中間那棵樹的果子，上帝曾說：『你們不可吃，也不可摸，免得你們死。』」
GEN|3|4|蛇對女人說：「你們不一定死；
GEN|3|5|因為上帝知道，你們吃的日子眼睛就開了，你們就像上帝一樣知道善惡。」
GEN|3|6|於是女人見那棵樹好作食物，又悅人的眼目，那樹令人喜愛，能使人有智慧，她就摘下果子吃了，又給了與她一起的丈夫，他也吃了。
GEN|3|7|他們二人的眼睛就開了，知道自己赤身露體，就編織無花果樹的葉子，為自己做成裙子。
GEN|3|8|天起了涼風，那人和他妻子聽見耶和華上帝在園中來回行走的聲音，就藏在園裏的樹木中，躲避耶和華上帝的面。
GEN|3|9|耶和華上帝呼喚那人，對他說：「你在哪裏？」
GEN|3|10|他說：「我在園中聽見你的聲音，我就害怕；因為我赤身露體，我就藏了起來。」
GEN|3|11|耶和華上帝說：「誰告訴你，你是赤身露體呢？莫非你吃了那樹上所出的，就是我吩咐你不可吃的嗎？」
GEN|3|12|那人說：「你賜給我、與我一起的女人，是她把那樹上所出的給我，我就吃了。」
GEN|3|13|耶和華上帝對女人說：「你怎麼會做這種事呢？」女人說：「那蛇引誘我，我就吃了。」
GEN|3|14|耶和華上帝對蛇說： 「你既做了這事，就必受詛咒， 比一切的牲畜和野獸更重。 你必用肚子行走， 終生吃土。
GEN|3|15|我要使你和女人彼此為仇， 你的後裔和女人的後裔也彼此為仇。 他要傷你的頭， 你要傷他的腳跟。 」
GEN|3|16|又對女人說： 「我必多多加增你懷胎的痛苦， 你生兒女時必多受痛苦。 你必戀慕你丈夫， 他必管轄你。」
GEN|3|17|又對 亞當 說： 「你既聽從你妻子的話， 吃了那樹上所出的， 就是我吩咐你不可吃的， 土地必因你的緣故受詛咒； 你必終生勞苦才能從土地得吃的。
GEN|3|18|土地必給你長出荊棘和蒺藜來； 你也要吃田間的五穀菜蔬。
GEN|3|19|你必汗流滿面才有食物可吃， 直到你歸了土地， 因為你是從土地而出的。 你本是塵土，仍要歸回塵土。」
GEN|3|20|那人給他妻子起名叫 夏娃 ，因為她是眾生之母 。
GEN|3|21|耶和華上帝用獸皮做衣服給 亞當 和他的妻子穿。
GEN|3|22|耶和華上帝說：「看哪，那人已經像我們中間的一個，知道善惡，現在恐怕他又伸手摘生命樹所出的來吃，就永遠活著。」
GEN|3|23|耶和華上帝就驅逐他出 伊甸園 ，使他耕種土地，他原是從土地裏被取出來的。
GEN|3|24|耶和華上帝把那人趕出去，就在 伊甸園 東邊安設基路伯和發出火焰轉動的劍，把守生命樹的道路。
GEN|4|1|那人和他妻子 夏娃 同房， 夏娃 就懷孕，生了 該隱 ，她說：「我靠耶和華得了一個男的。」
GEN|4|2|她又生了 該隱 的弟弟 亞伯 。 亞伯 是牧羊的； 該隱 是耕地的。
GEN|4|3|過了一些日子， 該隱 拿地裏的出產為供物獻給耶和華；
GEN|4|4|亞伯 也把他羊群中頭生的和羊的脂肪獻上。耶和華看中了 亞伯 和他的供物，
GEN|4|5|卻看不中 該隱 和他的供物。 該隱 就非常生氣，沉下臉來。
GEN|4|6|耶和華對 該隱 說：「你為甚麼生氣呢？你為甚麼沉下臉來呢？
GEN|4|7|你若做得對，豈不仰起頭來嗎？你若做得不對，罪就伏在門前。它想要控制你，你卻要制伏它。」
GEN|4|8|該隱 與他弟弟 亞伯 說話 。 二人正在田間時， 該隱 起來攻擊他弟弟 亞伯 ，把他殺了。
GEN|4|9|耶和華對 該隱 說：「你弟弟 亞伯 在哪裏？」他說：「我不知道！我豈是看守我弟弟的嗎？」
GEN|4|10|耶和華說：「你做了甚麼事呢？你弟弟血的聲音從地裏向我哀號。
GEN|4|11|現在你必從這地受詛咒，這地開了口，從你手裏接受你弟弟的血。
GEN|4|12|你耕種土地，它不再給你效力；你必流離飄蕩在地上。」
GEN|4|13|該隱 對耶和華說：「我的懲罰太重，過於我所能承當的。
GEN|4|14|看哪，今日你趕我離開這塊土地，不能見你的面；我必流離飄蕩在地上，凡遇見我的必殺我。」
GEN|4|15|耶和華對他說：「既然如此 ，凡殺 該隱 的，必遭報七倍。」耶和華就給 該隱 立一個記號，免得人遇見他就殺他。
GEN|4|16|於是 該隱 離開了耶和華的面，去住在 伊甸 東邊 挪得 之地。
GEN|4|17|該隱 與妻子同房，她就懷孕，生了 以諾 。 該隱 建造一座城，就照他兒子的名字稱那城為 以諾 。
GEN|4|18|以諾 生 以拿 ， 以拿 生 米戶雅利 ， 米戶雅利 生 瑪土撒利 ， 瑪土撒利 生 拉麥 。
GEN|4|19|拉麥 娶了兩個妻子：一個名叫 亞大 ，一個名叫 洗拉 。
GEN|4|20|亞大 生 雅八 ； 雅八 是住帳棚、牧養牲畜之人的祖師。
GEN|4|21|雅八 的兄弟名叫 猶八 ；他是所有彈琴吹簫之人的祖師。
GEN|4|22|洗拉 又生了 土八‧該隱 ；他是打造各樣銅器鐵器的工匠。 土八‧該隱 的妹妹是 拿瑪 。
GEN|4|23|拉麥 對他兩個妻子說： 亞大 、 洗拉 啊，聽我的聲音； 拉麥 的妻子啊，側耳聽我的言語： 大人傷我，我把他殺了； 小孩損我，我把他害了 。
GEN|4|24|若殺 該隱 ，遭報七倍， 殺 拉麥 的，必遭報七十七倍。
GEN|4|25|亞當 又與妻子同房，她就生了一個兒子，給他起名叫 塞特 ，說：「上帝給我立了另一個子嗣代替 亞伯 ，因為 該隱 殺了他。」
GEN|4|26|塞特 也生了一個兒子，起名叫 以挪士 。那時候，人開始求告耶和華的名。
GEN|5|1|這是 亞當 後代的家譜。當上帝造人的日子，他照著自己的樣式造人。
GEN|5|2|他造男造女。在他們被造的日子，上帝賜福給他們，稱他們為人。
GEN|5|3|亞當 活到一百三十歲，生了一個兒子，形像樣式和自己相似，就給他起名叫 塞特 。
GEN|5|4|亞當 生 塞特 之後，又活了八百年，並且生兒育女。
GEN|5|5|亞當 共活了九百三十年，就死了。
GEN|5|6|塞特 活到一百零五歲，生了 以挪士 。
GEN|5|7|塞特 生 以挪士 之後，又活了八百零七年，並且生兒育女。
GEN|5|8|塞特 共活了九百一十二年，就死了。
GEN|5|9|以挪士 活到九十歲，生了 該南 。
GEN|5|10|以挪士 生 該南 之後，又活了八百一十五年，並且生兒育女。
GEN|5|11|以挪士 共活了九百零五年，就死了。
GEN|5|12|該南 活到七十歲，生了 瑪勒列 。
GEN|5|13|該南 生 瑪勒列 之後，又活了八百四十年，並且生兒育女。
GEN|5|14|該南 共活了九百一十年，就死了。
GEN|5|15|瑪勒列 活到六十五歲，生了 雅列 。
GEN|5|16|瑪勒列 生 雅列 之後，又活了八百三十年，並且生兒育女。
GEN|5|17|瑪勒列 共活了八百九十五年，就死了。
GEN|5|18|雅列 活到一百六十二歲，生了 以諾 。
GEN|5|19|雅列 生 以諾 之後，又活了八百年，並且生兒育女。
GEN|5|20|雅列 共活了九百六十二年，就死了。
GEN|5|21|以諾 活到六十五歲，生了 瑪土撒拉 。
GEN|5|22|以諾 生 瑪土撒拉 之後，與上帝同行三百年，並且生兒育女。
GEN|5|23|以諾 共活了三百六十五年。
GEN|5|24|以諾 與上帝同行，上帝把他接去，他就不在了。
GEN|5|25|瑪土撒拉 活到一百八十七歲，生了 拉麥 。
GEN|5|26|瑪土撒拉 生 拉麥 之後，又活了七百八十二年，並且生兒育女。
GEN|5|27|瑪土撒拉 共活了九百六十九年，就死了。
GEN|5|28|拉麥 活到一百八十二歲，生了一個兒子，
GEN|5|29|給他起名叫 挪亞 ，說：「在耶和華所詛咒的地上，這個兒子必使我們從工作和手中的勞苦得到安慰。」
GEN|5|30|拉麥 生 挪亞 之後，又活了五百九十五年，並且生兒育女。
GEN|5|31|拉麥 共活了七百七十七年，就死了。
GEN|5|32|挪亞 活到五百歲，生了 閃 、 含 和 雅弗 。
GEN|6|1|當人開始在地面上增多、又生女兒的時候，
GEN|6|2|上帝的兒子們看見人的女子美貌，就隨意挑選，娶來為妻。
GEN|6|3|耶和華說：「人既屬乎血氣，我的靈就不永遠住在他裏面；然而他的年歲還可到一百二十年。」
GEN|6|4|那時候有巨人在地上，後來也有；上帝的兒子們和人的女子們交合，生了孩子。那些人就是古代的勇士，有名的人物。
GEN|6|5|耶和華見人在地上罪大惡極，終日心裏所想的盡都是惡事，
GEN|6|6|耶和華就因造人在地上感到遺憾，心中憂傷。
GEN|6|7|耶和華說：「我要把所造的人和走獸，爬行動物，以及天空的飛鳥，都從地面上除滅，因為我造了他們感到遺憾。」
GEN|6|8|只有 挪亞 在耶和華眼前蒙恩。
GEN|6|9|這是 挪亞 的後代。 挪亞 是個義人，在他的世代中是個完全人。 挪亞 與上帝同行。
GEN|6|10|挪亞 生了三個兒子，就是 閃 、 含 和 雅弗 。
GEN|6|11|這地在上帝面前敗壞了，地上充滿了暴力。
GEN|6|12|上帝觀看這地，看哪，它敗壞了，因為凡血肉之軀在地上的行為都敗壞了。
GEN|6|13|上帝對 挪亞 說：「在我面前，凡血肉之軀的結局已經臨到，因著他們，地上充滿了暴力。看哪，我要把他們和這地一起毀滅。
GEN|6|14|你要為自己用歌斐木造一艘方舟，並在方舟內造房間，內外都要抹上瀝青。
GEN|6|15|方舟的造法是這樣：要長三百肘，寬五十肘，高三十肘。
GEN|6|16|方舟上面要造天窗，向上一肘。方舟的門要開在旁邊。方舟要分上、中、下三層。
GEN|6|17|看哪，我要使洪水氾濫在地上，毀滅天下凡有生命氣息的血肉之軀，地上的一切都要滅亡。
GEN|6|18|但我要與你立約；你同你的兒子、妻子和媳婦都要進入方舟。
GEN|6|19|凡有血肉的動物，每樣一對，一公一母，你要帶進方舟，好跟你一起保全生命。
GEN|6|20|飛鳥各從其類，牲畜各從其類，地上的爬行動物各從其類，每樣一對，都要到你那裏，好保全生命。
GEN|6|21|你要拿各樣可吃的食物，儲存在你那裏，作你和牠們的糧食。」
GEN|6|22|挪亞 就去做了；凡上帝吩咐他的，他都照樣去做。
GEN|7|1|耶和華對 挪亞 說：「你和你的全家都要進入方舟，因為在這世代中，我看你在我面前是個義人。
GEN|7|2|凡潔淨的牲畜，你要各取七公七母；不潔淨的牲畜，你要各取一公一母；
GEN|7|3|天空的飛鳥也要各取七公七母，為了要留種，活在全地面上。
GEN|7|4|因為再過七天，我要降雨在地上四十晝夜，把我所造的一切生物從地面上除滅。」
GEN|7|5|挪亞 就遵照耶和華吩咐他的去做。
GEN|7|6|當洪水 在地上氾濫的時候， 挪亞 已六百歲。
GEN|7|7|挪亞 同他的兒子、妻子和媳婦都進入方舟，躲避洪水。
GEN|7|8|潔淨的牲畜和不潔淨的牲畜，飛鳥及所有爬行在土地上的，
GEN|7|9|都一對一對，有公有母，到 挪亞 那裏，進入方舟，正如上帝所吩咐 挪亞 的。
GEN|7|10|過了七天，洪水氾濫在地上。
GEN|7|11|挪亞 六百歲那一年的二月十七日，就在那一天，大深淵的泉源都裂開，天上的窗戶也敞開了，
GEN|7|12|四十晝夜有大雨降在地上。
GEN|7|13|正在那日， 挪亞 和他的兒子 閃 、 含 、 雅弗 ，以及 挪亞 的妻子和三個媳婦，都一同進入方舟。
GEN|7|14|他們和一切走獸，各從其類；一切牲畜，各從其類；地上爬的一切爬行動物，各從其類；一切的鳥，就是一切有翅膀的飛禽，各從其類；
GEN|7|15|凡有生命氣息的血肉之軀，都一對一對到 挪亞 那裏，進入方舟。
GEN|7|16|凡有血肉的，都一公一母進入方舟，正如上帝所吩咐 挪亞 的。耶和華就把他關在方舟裏。
GEN|7|17|洪水在地上氾濫四十天，水往上漲，使方舟浮起，方舟就從地上漂起來。
GEN|7|18|水勢洶湧，在地上大大上漲，方舟在水面上漂蕩。
GEN|7|19|水勢在地上極其浩大，普天下所有的高山都淹沒了。
GEN|7|20|水勢洶湧，比山高出十五肘 ，山嶺都淹沒了。
GEN|7|21|凡有血肉在地上行動的，就是飛鳥、牲畜、走獸和地上成群的群聚動物，以及所有的人，都死了。
GEN|7|22|在乾地上凡鼻孔裏有生命氣息的都死了。
GEN|7|23|耶和華除滅了地面上各類的生物，包括人和牲畜、爬行動物，以及天空的飛鳥；他們就都從地上除滅了，只剩下 挪亞 和那些與他同在方舟裏的。
GEN|7|24|水勢洶湧，在地上共一百五十天。
GEN|8|1|上帝記念 挪亞 和 挪亞 方舟裏的一切走獸牲畜。上帝使風吹地，水勢漸落。
GEN|8|2|深淵的泉源和天上的窗戶都關閉了，雨不再從天降下。
GEN|8|3|水從地上逐漸消退。過了一百五十天，水就退了。
GEN|8|4|七月十七日，方舟停在 亞拉臘山 上。
GEN|8|5|水繼續退去，直到十月；十月初一，山頂都露出來了。
GEN|8|6|過了四十天， 挪亞 打開他所造的方舟的窗戶，
GEN|8|7|放出一隻烏鴉。那烏鴉飛來飛去，直到地上的水都乾了。
GEN|8|8|他又從他那裏放出一隻鴿子，要看水從地面上退了沒有。
GEN|8|9|但全地面都是水，鴿子找不到落腳之地，就回到方舟 挪亞 那裏。 挪亞 伸手接了鴿子，把牠帶進方舟。
GEN|8|10|挪亞 又另外等了七天，再把鴿子從方舟放出去。
GEN|8|11|到了晚上，鴿子回到他那裏，看哪，嘴裏有一片剛啄下來的橄欖葉， 挪亞 就知道水已經從地上退了。
GEN|8|12|他又另外等了七天，再放出鴿子，這次鴿子不再回到他那裏了。
GEN|8|13|當 挪亞 六百零一歲，正月初一的時候，地上的水都乾了。 挪亞 打開方舟的蓋觀看，看哪，地面乾了。
GEN|8|14|到了二月二十七日，地就都乾了。
GEN|8|15|上帝對 挪亞 說：
GEN|8|16|「你同你的妻子、兒子、媳婦都要出方舟。
GEN|8|17|凡與你一起有血肉的生物，就是飛鳥、牲畜和地上爬的一切爬行動物，都要帶出來。 牠們要在地上滋生，繁殖增多。」
GEN|8|18|於是 挪亞 同他的兒子、妻子、媳婦都出來了。
GEN|8|19|一切走獸、爬行動物和飛鳥，地上所有的動物，各從其類，也都出了方舟。
GEN|8|20|挪亞 為耶和華築了一座壇，拿各種潔淨的牲畜和各種潔淨的飛鳥，獻在壇上為燔祭。
GEN|8|21|耶和華聞了那馨香之氣，耶和華心裏說：「我不再因人的緣故詛咒土地，因為人從幼年就心裏懷著惡念；我也不再照我曾做的毀滅一切生物了。
GEN|8|22|地還存在的時候，撒種、收割、寒暑、冬夏、晝夜都永不止息。」
GEN|9|1|上帝賜福給 挪亞 和他的兒子，對他們說：「你們要生養眾多，遍滿這地。
GEN|9|2|地上一切的走獸、天空一切的飛鳥、所有爬行在土地上的和海裏一切的魚都必怕你們，畏懼你們，牠們都要交在你們手裏。
GEN|9|3|凡活的動物都可作你們的食物。這一切我都賜給你們，如同綠色的菜蔬一樣。
GEN|9|4|只是帶著生命的肉，就是帶著血的，你們不可吃。
GEN|9|5|流你們血、害你們命的，我必向他追討；我要向一切走獸追討，向人和向人的弟兄追討人命。
GEN|9|6|凡流人血的，他的血也必被人所流，因為上帝造人，是照自己的形像造的。
GEN|9|7|你們要生養眾多，在地上繁衍昌盛。」
GEN|9|8|上帝對 挪亞 和同他一起的兒子說：
GEN|9|9|「看哪，我要與你們和你們後裔立我的約，
GEN|9|10|包括和你們一起所有的生物，就是飛鳥、牲畜、地上一切的走獸，凡從方舟裏出來地上一切的生物。
GEN|9|11|我與你們立我的約：凡有血肉的，不再被洪水滅絕，也不再有洪水毀壞這地了。」
GEN|9|12|上帝說：「這是我與你們，以及和你們一起的一切生物所立之約的記號，直到萬代：
GEN|9|13|我把彩虹放在雲中，這就是我與地立約的記號了。
GEN|9|14|我使雲遮地的時候，會有彩虹出現在雲中，
GEN|9|15|我就記念我與你們，以及各樣有血肉的生物所立的約：不再有洪水氾濫去毀滅一切有血肉的了。
GEN|9|16|彩虹出現在雲中，我看見了，就要記念上帝與地上一切有血肉的生物所立的永約。」
GEN|9|17|上帝對 挪亞 說：「這就是我與地上一切有血肉的立約的記號。」
GEN|9|18|挪亞 的兒子，從方舟出來的，有 閃 、 含 和 雅弗 。 含 是 迦南 的父親。
GEN|9|19|這是 挪亞 的三個兒子，他們的後裔散佈全地。
GEN|9|20|挪亞 是農夫，是他開始栽葡萄園的。
GEN|9|21|他喝了一些酒就醉了，在他的帳棚裏赤著身子。
GEN|9|22|迦南 的父親 含 看見他父親赤身，就到外面告訴他的兩個兄弟。
GEN|9|23|於是 閃 和 雅弗 拿了外衣搭在二人肩上，倒退著進去，遮蓋父親的赤身；他們背著臉，看不見父親的赤身。
GEN|9|24|挪亞 酒醒以後，知道小兒子向他所做的事，
GEN|9|25|就說： 「 迦南 當受詛咒， 必給他弟兄作奴僕的奴僕。」
GEN|9|26|又說： 「耶和華— 閃 的上帝是應當稱頌的！ 願 迦南 作 閃 的奴僕。
GEN|9|27|願上帝使 雅弗 擴張， 願他住在 閃 的帳棚裏； 願 迦南 作他的奴僕。」
GEN|9|28|洪水以後， 挪亞 又活了三百五十年。
GEN|9|29|挪亞 共活了九百五十年，就死了。
GEN|10|1|這是 挪亞 的兒子 閃 、 含 、 雅弗 的後代。洪水以後，他們都生了兒子。
GEN|10|2|雅弗 的兒子是 歌篾 、 瑪各 、 瑪代 、 雅完 、 土巴 、 米設 、 提拉 。
GEN|10|3|歌篾 的兒子是 亞實基拿 、 利法 、 陀迦瑪 。
GEN|10|4|雅完 的兒子是 以利沙 、 他施 、 基提 、 羅單 人 。
GEN|10|5|從這些人中有沿海國家的人散居各處，有自己的土地，各有各的語言、宗族、國家。
GEN|10|6|含 的兒子是 古實 、 麥西 、 弗 、 迦南 。
GEN|10|7|古實 的兒子是 西巴 、 哈腓拉 、 撒弗他 、 拉瑪 、 撒弗提迦 。 拉瑪 的兒子是 示巴 、 底但 。
GEN|10|8|古實 又生 寧錄 ，他是地上第一個勇士。
GEN|10|9|他在耶和華面前是個英勇的獵人，所以有話說：「像 寧錄 在耶和華面前是個英勇的獵人。」
GEN|10|10|他王國的開始是在 巴別 、 以力 、 亞甲 、 甲尼 ，都在 示拿 地。
GEN|10|11|他從那地出來往 亞述 去，建造了 尼尼微 、 利河伯 、 迦拉 ，
GEN|10|12|以及 尼尼微 和 迦拉 之間的 利鮮 ，那是座大城。
GEN|10|13|麥西 生 路低 人、 亞拿米 人、 利哈比 人、 拿弗土希 人、
GEN|10|14|帕斯魯細 人、 迦斯路希 人、 迦斐託 人； 非利士 人是從 迦斐託 人 出來的。
GEN|10|15|迦南 生了長子 西頓 ，又生 赫
GEN|10|16|和 耶布斯 人、 亞摩利 人、 革迦撒 人、
GEN|10|17|希未 人、 亞基 人、 西尼 人、
GEN|10|18|亞瓦底 人、 洗瑪利 人、 哈馬 人，後來 迦南 的家族散開了。
GEN|10|19|迦南 的疆界是從 西頓 到 基拉耳 ，直到 迦薩 ，又到 所多瑪 、 蛾摩拉 、 押瑪 、 洗扁 ，直到 拉沙 。
GEN|10|20|這就是 含 的後裔，各有自己的宗族、語言、土地和國家。
GEN|10|21|閃 也生了兒子，他是 雅弗 的哥哥 ，是 希伯 人的祖先。
GEN|10|22|閃 的兒子是 以攔 、 亞述 、 亞法撒 、 路德 、 亞蘭 。
GEN|10|23|亞蘭 的兒子是 烏斯 、 戶勒 、 基帖 、 瑪施 。
GEN|10|24|亞法撒 生 沙拉 ， 沙拉 生 希伯 。
GEN|10|25|希伯 生了兩個兒子，一個名叫 法勒 ，因為那時人分地居住； 法勒 的兄弟名叫 約坍 。
GEN|10|26|約坍 生 亞摩答 、 沙列 、 哈薩瑪非 、 耶拉 、
GEN|10|27|哈多蘭 、 烏薩 、 德拉 、
GEN|10|28|俄巴路 、 亞比瑪利 、 示巴 、
GEN|10|29|阿斐 、 哈腓拉 、 約巴 ，這些都是 約坍 的兒子。
GEN|10|30|他們所住的地方是從 米沙 直到 西發 ，到東邊的山。
GEN|10|31|這就是 閃 的後裔，各有自己的宗族、語言、土地和國家。
GEN|10|32|這些是 挪亞 兒子的宗族，按著他們的後代立國。洪水以後，邦國就從他們散佈在地上。
GEN|11|1|那時，全地只有一種語言，都說一樣的話。
GEN|11|2|他們向東遷移的時候，在 示拿 地找到一片平原，就住在那裏。
GEN|11|3|他們彼此商量說：「來，讓我們來做磚，把磚燒透了。」他們就拿磚當石頭，又拿柏油當泥漿。
GEN|11|4|他們說：「來，讓我們建造一座城和一座塔，塔頂通天。我們要為自己立名，免得我們分散在全地面上。」
GEN|11|5|耶和華降臨，要看世人所建造的城和塔。
GEN|11|6|耶和華說：「看哪，他們成了同一個民族，都有一樣的語言。這只是他們開始做的事，現在他們想要做的任何事，就沒有甚麼可攔阻他們了。
GEN|11|7|來，我們下去，在那裏變亂他們的語言，使他們彼此語言不通。」
GEN|11|8|於是耶和華使他們從那裏分散在全地面上；他們就停止建造那城了。
GEN|11|9|因為耶和華在那裏變亂了全地的語言，把人從那裏分散在全地面上，所以那城名叫 巴別 。
GEN|11|10|這是 閃 的後代。洪水以後二年， 閃 一百歲生了 亞法撒 。
GEN|11|11|閃 生 亞法撒 之後又活了五百年，並且生兒育女。
GEN|11|12|亞法撒 活到三十五歲，生了 沙拉 。
GEN|11|13|亞法撒 生 沙拉 之後又活了四百零三年，並且生兒育女。
GEN|11|14|沙拉 活到三十歲，生了 希伯 。
GEN|11|15|沙拉 生 希伯 之後又活了四百零三年，並且生兒育女。
GEN|11|16|希伯 活到三十四歲，生了 法勒 。
GEN|11|17|希伯 生 法勒 之後又活了四百三十年，並且生兒育女。
GEN|11|18|法勒 活到三十歲，生了 拉吳 。
GEN|11|19|法勒 生 拉吳 之後又活了二百零九年，並且生兒育女。
GEN|11|20|拉吳 活到三十二歲，生了 西鹿 。
GEN|11|21|拉吳 生 西鹿 之後又活了二百零七年，並且生兒育女。
GEN|11|22|西鹿 活到三十歲，生了 拿鶴 。
GEN|11|23|西鹿 生 拿鶴 之後又活了二百年，並且生兒育女。
GEN|11|24|拿鶴 活到二十九歲，生了 他拉 。
GEN|11|25|拿鶴 生 他拉 之後又活了一百一十九年，並且生兒育女。
GEN|11|26|他拉 活到七十歲，生了 亞伯蘭 、 拿鶴 和 哈蘭 。
GEN|11|27|這是 他拉 的後代。 他拉 生 亞伯蘭 、 拿鶴 和 哈蘭 ； 哈蘭 生 羅得 。
GEN|11|28|哈蘭 死在他父親 他拉 的面前，死在他的出生地 迦勒底 的 吾珥 。
GEN|11|29|亞伯蘭 、 拿鶴 各娶了妻。 亞伯蘭 的妻子名叫 撒萊 ， 拿鶴 的妻子名叫 密迦 ，是 哈蘭 的女兒。 哈蘭 是 密迦 和 亦迦 的父親。
GEN|11|30|撒萊 不生育，沒有孩子。
GEN|11|31|他拉 帶著他兒子 亞伯蘭 和他孫子， 哈蘭 的兒子 羅得 ，以及他的媳婦， 亞伯蘭 的妻子 撒萊 ，一同出了 迦勒底 的 吾珥 ，要往 迦南 地去；他們來到 哈蘭 ，就住在那裏。
GEN|11|32|他拉 共活了二百零五年，就死在 哈蘭 。
GEN|12|1|耶和華對 亞伯蘭 說：「你要離開本地、本族、父家，往我所要指示你的地去。
GEN|12|2|我必使你成為大國，我必賜福給你，使你的名為大；你要使別人得福 。
GEN|12|3|為你祝福的，我必賜福給他；詛咒你的，我必詛咒他。地上的萬族都必因你得福。」
GEN|12|4|亞伯蘭 就遵照耶和華的吩咐去了； 羅得 也和他同去。 亞伯蘭 離開 哈蘭 的時候年七十五歲。
GEN|12|5|亞伯蘭 帶著他妻子 撒萊 和姪兒 羅得 ，以及他們在 哈蘭 積蓄的財物、獲得的人口，往 迦南 地去。他們就來到了 迦南 地。
GEN|12|6|亞伯蘭 經過那地，直到 示劍 地方， 摩利 橡樹那裏；當時 迦南 人住在那地。
GEN|12|7|耶和華向 亞伯蘭 顯現，說：「我要把這地賜給你的後裔。」 亞伯蘭 就在那裏為向他顯現的耶和華築了一座壇。
GEN|12|8|從那裏他又遷到 伯特利 東邊的山，支搭帳棚；西邊是 伯特利 ，東邊是 艾 。他在那裏又為耶和華築了一座壇，求告耶和華的名。
GEN|12|9|後來 亞伯蘭 漸漸遷往 尼革夫 去。
GEN|12|10|那地遭遇饑荒。 亞伯蘭 因那地的饑荒嚴重，就下到 埃及 ，要在那裏寄居。
GEN|12|11|將近 埃及 ，他對妻子 撒萊 說：「看哪，我知道你是美貌的女人。
GEN|12|12|埃及 人看見你會說：『這是他的妻子』，他們就會殺我，卻讓你活著。
GEN|12|13|所以，請你說你是我的妹妹，使我可以因你得平安，我的性命也因你存活。」
GEN|12|14|亞伯蘭 到達 埃及 時， 埃及 人看見那女人極其美貌。
GEN|12|15|法老的臣僕看見了她，就在法老面前稱讚她。那女人就被帶進法老的宮中。
GEN|12|16|法老就因她厚待 亞伯蘭 ，給了 亞伯蘭 許多牛、羊、公驢、奴僕、婢女、母驢、駱駝。
GEN|12|17|耶和華因 亞伯蘭 妻子 撒萊 的緣故，降大災擊打法老和他的全家。
GEN|12|18|法老召了 亞伯蘭 來，說：「你向我做的是甚麼事呢？為甚麼沒有告訴我她是你的妻子？
GEN|12|19|為甚麼說『她是我的妹妹』，以致我把她接來要作我的妻子呢？現在 ，看哪，你的妻子在這裏，帶她走吧！」
GEN|12|20|於是法老吩咐人把 亞伯蘭 和他妻子，以及他一切所有的都送走了。
GEN|13|1|亞伯蘭 帶著他的妻子與 羅得 ，以及一切所有的，從 埃及 上 尼革夫 去。
GEN|13|2|亞伯蘭 的牲畜和金銀極多。
GEN|13|3|他從 尼革夫 漸漸往 伯特利 去，到了 伯特利 和 艾 的中間，當初他支搭帳棚的地方，
GEN|13|4|也是他起先築壇的地方。 亞伯蘭 在那裏求告耶和華的名。
GEN|13|5|與 亞伯蘭 同行的 羅得 也有牛群、羊群、帳棚。
GEN|13|6|那地容不下他們住在一起；因為他們的財物非常多，使他們不能同住一起。
GEN|13|7|當時， 迦南 人與 比利洗 人在那地居住。 亞伯蘭 的牧人和 羅得 的牧人之間起了爭端。
GEN|13|8|亞伯蘭 就對 羅得 說：「你我不可以相爭，你的牧人和我的牧人也不可以相爭，因為我們是一家人。
GEN|13|9|遍地不都在你眼前嗎？請你離開我吧！你向左，我就向右；你向右，我就向左。」
GEN|13|10|羅得 舉目，看見 約旦河 整個平原，直到 瑣珥 ，都是水源充足之地。在耶和華未毀滅 所多瑪 、 蛾摩拉 以前，那地好像耶和華的園子，又像 埃及 地。
GEN|13|11|於是 羅得 選擇了 約旦河 整個平原。 羅得 往東遷移，他們就彼此分開了。
GEN|13|12|亞伯蘭 住在 迦南 地； 羅得 住在平原的城鎮，他漸漸遷移帳棚，直到 所多瑪 。
GEN|13|13|所多瑪 人在耶和華面前罪大惡極。
GEN|13|14|羅得 離開 亞伯蘭 以後，耶和華對 亞伯蘭 說：「你要從你所在的地方，舉目向東西南北觀看；
GEN|13|15|你所看見一切的地，我都要把它賜給你和你的後裔，直到永遠。
GEN|13|16|我要使你的後裔好像地上的塵沙，人若能數地上的塵沙，才能數你的後裔。
GEN|13|17|你起來，縱橫走遍這地，因為我必把這地賜給你。」
GEN|13|18|亞伯蘭 就遷移帳棚，來到 希伯崙 ， 幔利 的橡樹那裏居住，在那裏為耶和華築了一座壇。
GEN|14|1|當 暗拉非 作 示拿 王， 亞略 作 以拉撒 王， 基大老瑪 作 以攔 王， 提達 作 戈印 王的時候，
GEN|14|2|他們攻打 所多瑪 王 比拉 、 蛾摩拉 王 比沙 、 押瑪 王 示納 、 洗扁 王 善以別 和 比拉 王， 比拉 就是 瑣珥 。
GEN|14|3|這些王都會合在 西訂谷 ， 西訂谷 就是 鹽海 。
GEN|14|4|他們已經服事 基大老瑪 十二年，第十三年就背叛了。
GEN|14|5|第十四年， 基大老瑪 和與他結盟的王都來了，在 亞特律‧加寧 擊敗 利乏音 人，在 哈麥 擊敗 蘇西 人，在 沙微‧基列亭 擊敗 以米 人，
GEN|14|6|在 何利 人的 西珥山 擊敗 何利 人，一直到靠近曠野的 伊勒‧巴蘭 。
GEN|14|7|他們轉回，來到 安‧密巴 ，就是 加低斯 ，擊敗了 亞瑪力 全地的人，以及住在 哈洗遜‧他瑪 的 亞摩利 人。
GEN|14|8|於是 所多瑪 王、 蛾摩拉 王、 押瑪 王、 洗扁 王和 比拉 王， 比拉 就是 瑣珥 ，都出來，在 西訂谷 擺陣，與他們交戰，
GEN|14|9|就是與 以攔 王 基大老瑪 、 戈印 王 提達 、 示拿 王 暗拉非 、 以拉撒 王 亞略 交戰；這就是四王對五王之戰。
GEN|14|10|西訂谷 有許多柏油坑。 所多瑪 王和 蛾摩拉 王逃跑，掉在坑裏，其餘的人都往山上逃跑。
GEN|14|11|四王就把 所多瑪 和 蛾摩拉 所有的財物和所有的糧食都擄掠去了；
GEN|14|12|他們也把 亞伯蘭 的姪兒 羅得 和 羅得 的財物都擄掠去了。當時 羅得 住在 所多瑪 。
GEN|14|13|有一個逃脫的人來告訴 希伯來 人 亞伯蘭 ； 亞伯蘭 正住在 亞摩利 人 幔利 的橡樹那裏。 幔利 、 以實各 和 亞乃 都是弟兄，曾與 亞伯蘭 結盟。
GEN|14|14|亞伯蘭 聽見他姪兒 被擄去，就把三百一十八個生在他家中、受過訓練的壯丁全都出動 去追，一直到 但 。
GEN|14|15|在夜間，他和他的僕人分隊擊敗了敵人，並且追殺他們，直到 大馬士革 北邊的 何把 。
GEN|14|16|他把一切被擄掠的財物奪回，也把他姪兒 羅得 和他的財物，以及人和婦女都奪回來。
GEN|14|17|亞伯蘭 擊敗 基大老瑪 和與他結盟的王回來的時候， 所多瑪 王出來，在 沙微谷 迎接他， 沙微谷 就是 王的谷 。
GEN|14|18|又有 撒冷 王 麥基洗德 帶著餅和酒出來；他是至高上帝的祭司。
GEN|14|19|他為 亞伯蘭 祝福，說： 「願至高的上帝、 天地的主賜福給 亞伯蘭 ！
GEN|14|20|至高的上帝把敵人交在你手裏， 他是應當稱頌的！」 亞伯蘭 就把所有的拿出十分之一給他。
GEN|14|21|所多瑪 王對 亞伯蘭 說：「你把人還給我，財物你自己拿去吧！」
GEN|14|22|亞伯蘭 對 所多瑪 王說：「我指著耶和華—至高的上帝、天地的主起誓：
GEN|14|23|凡是你的東西，就是一根線、一條鞋帶，我都不拿，免得你說：『是我使 亞伯蘭 富足！』
GEN|14|24|我甚麼都不要，只是僕人所吃的，以及與我同去的 亞乃 、 以實各 、 幔利 所應得的份，讓他們拿去吧！」
GEN|15|1|這些事以後，耶和華的話在異象中臨到 亞伯蘭 ，說：「 亞伯蘭 哪，不要懼怕！我是你的盾牌，你必得豐富的賞賜。」
GEN|15|2|亞伯蘭 說：「主耶和華啊，我還沒有兒子，你能賜我甚麼呢？承受我家業的是 大馬士革 人 以利以謝 。」
GEN|15|3|亞伯蘭 又說：「看哪，你沒有給我後嗣。你看，那生在我家中的人要繼承我。」
GEN|15|4|看哪，耶和華的話又臨到他，說：「這人不會繼承你，你本身所生的才會繼承你。」
GEN|15|5|於是耶和華帶他到外面，說：「你向天觀看，去數星星，你能數得清嗎？」又對他說：「你的後裔將要如此。」
GEN|15|6|亞伯蘭 信耶和華，耶和華就以此算他為義。
GEN|15|7|耶和華又對他說：「我是耶和華，曾領你出 迦勒底 的 吾珥 ，為要把這地賜你為業。」
GEN|15|8|亞伯蘭 說：「主耶和華啊，我怎能知道我必得這地為業呢？」
GEN|15|9|耶和華對他說：「你為我取一頭三歲的母牛犢，一隻三歲的母山羊，一隻三歲的公綿羊，一隻斑鳩和一隻雛鴿。」
GEN|15|10|亞伯蘭 就把這些都取來，每樣從中間劈成兩半，一半對著另一半排列，只有鳥沒有劈開。
GEN|15|11|當鷙鳥下來，落在這些屍體上時， 亞伯蘭 就把牠們趕走了。
GEN|15|12|日落的時候， 亞伯蘭 沉睡了。看哪，有大而可怕的黑暗落在他身上。
GEN|15|13|耶和華對 亞伯蘭 說：「你要確實知道，你的後裔必寄居在別人的地，服事那地的人；那地的人要虐待他們四百年。
GEN|15|14|但我要懲罰他們所服事的那國，以後他們必帶著許多財物從那裏出來。
GEN|15|15|至於你，你要平平安安歸到你祖先那裏，必享長壽，被人埋葬。
GEN|15|16|到了第四代，他們必回到這裏，因為 亞摩利 人的罪惡到現在還沒有滿盈。」
GEN|15|17|日落天黑的時候，看哪，有冒煙的爐和燒著的火把從那些肉塊中經過。
GEN|15|18|在那日，耶和華與 亞伯蘭 立約，說：「我已賜給你的後裔這一片地，從 埃及河 直到 大河 ， 幼發拉底河 ，
GEN|15|19|就是 基尼 人、 基尼洗 人、 甲摩尼 人、
GEN|15|20|赫 人、 比利洗 人、 利乏音 人、
GEN|15|21|亞摩利 人、 迦南 人、 革迦撒 人、 耶布斯 人的地。」
GEN|16|1|亞伯蘭 的妻子 撒萊 沒有為他生孩子。 撒萊 有一個婢女，是 埃及 人，名叫 夏甲 。
GEN|16|2|撒萊 對 亞伯蘭 說：「看哪，耶和華使我不能生育。你來和我的婢女同房，也許我可以從她得孩子 。」 亞伯蘭 聽從了 撒萊 的話。
GEN|16|3|於是 亞伯蘭 的妻子 撒萊 把她的婢女， 埃及 人 夏甲 ，給了丈夫為妾；那時 亞伯蘭 在 迦南 已經住了十年。
GEN|16|4|亞伯蘭 與 夏甲 同房， 夏甲 就懷了孕。她看見自己有孕，就輕視她的女主人。
GEN|16|5|撒萊 對 亞伯蘭 說：「我因你受了委屈。我把我的婢女放在你懷中，她見自己懷了孕，就輕視我。願耶和華在你我之間判斷。」
GEN|16|6|亞伯蘭 對 撒萊 說：「看哪，婢女在你手裏，你可以照你看為好的對待她。」於是， 撒萊 虐待她，她就從 撒萊 面前逃走了。
GEN|16|7|耶和華的使者在曠野的水泉旁，在 書珥 路上的水泉旁遇見 夏甲 ，
GEN|16|8|對她說：「 撒萊 的婢女 夏甲 ，你從哪裏來？要到哪裏去？」她說：「我從我的女主人 撒萊 面前逃出來。」
GEN|16|9|耶和華的使者對她說：「你要回到你的女主人那裏，屈服在她手下。」
GEN|16|10|耶和華的使者對她說： 「我必使你的後裔極其繁多， 多到不可勝數。」
GEN|16|11|耶和華的使者又對她說： 「看哪，你已懷孕， 要生一個兒子。 你要給他起名叫 以實瑪利 ， 因為耶和華聽見了你的苦楚。
GEN|16|12|他為人必像野驢。 他的手要攻打人， 人的手也要攻打他； 他必常與他的眾弟兄作對 。」
GEN|16|13|夏甲 就稱那向她說話的耶和華為「你是看見 的上帝」，因為她說：「他看見了我之後，我還能在這裏看見他嗎？」
GEN|16|14|所以這井名叫 庇耳‧拉海‧萊 ，看哪，它位於 加低斯 和 巴列 的中間。
GEN|16|15|後來 夏甲 為 亞伯蘭 生了一個兒子； 亞伯蘭 給 夏甲 生的兒子起名叫 以實瑪利 。
GEN|16|16|夏甲 為 亞伯蘭 生 以實瑪利 的時候， 亞伯蘭 年八十六歲。
GEN|17|1|亞伯蘭 九十九歲時，耶和華向他顯現，對他說：「我是全能的上帝。你當在我面前行走，作完全的人，
GEN|17|2|我要與你立約，使你的後裔極其繁多。」
GEN|17|3|亞伯蘭 臉伏於地；上帝又對他說：
GEN|17|4|「看哪，這就是我與你立的約，你要成為多國的父。
GEN|17|5|從今以後，你的名字不再叫 亞伯蘭 ，要叫 亞伯拉罕 ，因為我已經立你作多國之父。
GEN|17|6|我必使你生養極其繁多；國度要從你而立，君王要從你而出。
GEN|17|7|我要與你，以及你世世代代的後裔堅立我的約，成為永遠的約，是要作你和你後裔的上帝。
GEN|17|8|我要把你現在寄居的地，就是 迦南 全地，賜給你和你的後裔永遠為業；我也必作他們的上帝。」
GEN|17|9|上帝又對 亞伯拉罕 說：「你和你的後裔一定要世世代代遵守我的約。
GEN|17|10|這就是我與你，以及你的後裔所立的約，是你們所當遵守的，你們所有的男子都要受割禮。
GEN|17|11|你們要割去肉體的包皮，這是我與你們立約的記號。
GEN|17|12|你們世世代代的男子，無論是在家裏生的，或是用銀子從外人買來而不是你後裔生的，都要在生下來的第八日受割禮。
GEN|17|13|你家裏生的和你用銀子買的，都必須受割禮。這樣，我的約就在你們肉體上成為永遠的約。
GEN|17|14|不受割禮的男子都必從民中剪除，因他違背了我的約。」
GEN|17|15|上帝又對 亞伯拉罕 說：「至於你的妻子 撒萊 ，不可再叫她 撒萊 ，她的名要叫 撒拉 。
GEN|17|16|我必賜福給她，也要從她賜一個兒子給你。我必賜福給 撒拉 ，她要興起多國；必有百姓的君王從她而出。」
GEN|17|17|亞伯拉罕 就臉伏於地竊笑，心裏想：「一百歲的人還能有孩子嗎？ 撒拉 已經九十歲了，還能生育嗎？」
GEN|17|18|亞伯拉罕 對上帝說：「但願 以實瑪利 活在你面前。」
GEN|17|19|上帝說：「不！你妻子 撒拉 必為你生一個兒子，你要給他起名叫 以撒 。我要與他堅立我的約，成為他後裔永遠的約。
GEN|17|20|至於 以實瑪利 ，我已聽見你了：看哪，我必賜福給他，使他興旺，極其繁多。他必生十二個族長，我要使他成為大國。
GEN|17|21|到明年所定的時候， 撒拉 必為你生 以撒 ，我要與他堅立我的約。」
GEN|17|22|上帝和 亞伯拉罕 說完了話，就離開他上升去了。
GEN|17|23|在那一天， 亞伯拉罕 遵照上帝所說的，給他的兒子 以實瑪利 和家裏所有的男丁，無論是在家裏生的，或是用銀子買來的，都行了割禮 。
GEN|17|24|亞伯拉罕 受割禮時，年九十九歲。
GEN|17|25|他兒子 以實瑪利 受割禮時，年十三歲。
GEN|17|26|在那一天， 亞伯拉罕 和他兒子 以實瑪利 一同受了割禮。
GEN|17|27|家裏所有的男人，無論是在家裏生的，或是用銀子從外人買來的，也都一同受了割禮。
GEN|18|1|耶和華在 幔利 橡樹那裏向 亞伯拉罕 顯現。天正熱的時候， 亞伯拉罕 坐在帳棚門口。
GEN|18|2|他舉目觀看，看哪，有三個人站在他附近。他一看見，就從帳棚門口跑去迎接他們，俯伏在地，
GEN|18|3|說：「我主，我若在你眼前蒙恩，請不要離開你的僕人走過去。
GEN|18|4|容我拿點水來，請你們洗腳，在樹下休息。
GEN|18|5|既然你們來到僕人這裏了，我再拿點餅來，讓你們恢復心力，然後再走。」他們說：「就照你說的去做吧。」
GEN|18|6|亞伯拉罕 急忙進帳棚到 撒拉 那裏，說：「你趕快拿三細亞細麵，揉麵做餅。」
GEN|18|7|亞伯拉罕 又跑到牛群裏，牽了一頭又嫩又好的牛犢來，交給僕人，僕人就急忙去預備。
GEN|18|8|亞伯拉罕 取了乳酪和奶，以及預備好了的牛犢來，擺在他們面前，自己在樹下站在旁邊，他們就吃了。
GEN|18|9|他們對 亞伯拉罕 說：「你妻子 撒拉 在哪裏？」他說：「看哪，在帳棚裏。」
GEN|18|10|有一位說：「明年這時候 ，我一定會回到你這裏。看哪，你的妻子 撒拉 會生一個兒子。」 撒拉 在那人後面的帳棚門口也聽見了。
GEN|18|11|亞伯拉罕 和 撒拉 都年紀老邁， 撒拉 的月經已停了。
GEN|18|12|撒拉 心裏竊笑，說：「我已衰老，我的主也老了，怎能有這喜事呢？」
GEN|18|13|耶和華對 亞伯拉罕 說：「 撒拉 為甚麼竊笑，說：『我已年老，果真能生育嗎？』
GEN|18|14|耶和華豈有難成的事嗎？到了所定的時候，我必回到你這裏。明年這時候， 撒拉 會生一個兒子。」
GEN|18|15|撒拉 因為害怕，就不承認，說：「我沒有笑。」那人說：「不，你的確笑了。」
GEN|18|16|三人從那裏起程，面向 所多瑪 觀望， 亞伯拉罕 與他們同行，要送他們一程。
GEN|18|17|耶和華說：「我所要做的事豈可瞞著 亞伯拉罕 呢？
GEN|18|18|亞伯拉罕 必要成為強大的國；地上的萬國都必因他得福。
GEN|18|19|我揀選他 ，為要叫他命令他的子孫和後代家屬遵行耶和華的道，秉公行義，使耶和華所應許 亞伯拉罕 的話都實現了。」
GEN|18|20|耶和華說：「 所多瑪 和 蛾摩拉 罪惡極其嚴重，控告他們的聲音很大。
GEN|18|21|我要下去察看他們所做的，是否真的像那達到我這裏的聲音一樣；如果不是，我也要知道。」
GEN|18|22|二人轉身離開那裏，往 所多瑪 去；但 亞伯拉罕 仍然站在耶和華面前。
GEN|18|23|亞伯拉罕 近前來，說：「你真的要把義人和惡人一同剿滅嗎？
GEN|18|24|假若那城裏有五十個義人，你真的還要剿滅，不因城裏這五十個義人饒了那地方嗎？
GEN|18|25|你絕不會做這樣的事，把義人與惡人一同殺了，使義人與惡人一樣。你絕不會這樣！審判全地的主豈不做公平的事嗎？」
GEN|18|26|耶和華說：「我若在 所多瑪城 裏找到五十個義人，我就為他們的緣故饒恕那整個地方。」
GEN|18|27|亞伯拉罕 回答說：「看哪，我雖只是塵土灰燼，還敢向主說話。
GEN|18|28|假若這五十個義人少了五個，你就因為少了五個而毀滅全城嗎？」他說：「我在那裏若找到四十五個，就不毀滅。」
GEN|18|29|亞伯拉罕 又對他說：「假若在那裏找到四十個呢？」他說：「為這四十個的緣故，我也不做。」
GEN|18|30|亞伯拉罕 說：「求主不要生氣，容我說，假若在那裏找到三十個呢？」他說：「我在那裏若找到三十個，我也不做。」
GEN|18|31|亞伯拉罕 說：「看哪，我還敢向主說，假若在那裏找到二十個呢？」他說：「為這二十個的緣故，我也不毀滅。」
GEN|18|32|亞伯拉罕 說：「求主不要生氣，我再說一次，假若在那裏找到十個呢？」他說：「為這十個的緣故，我也不毀滅。」
GEN|18|33|耶和華與 亞伯拉罕 說完了話就走了； 亞伯拉罕 也回到自己的地方去了。
GEN|19|1|兩個天使在傍晚到了 所多瑪 ， 羅得 正坐在 所多瑪 的城門口。 羅得 一看見，就起身迎接他們，臉伏於地下拜，
GEN|19|2|說：「看哪，我主，請你們轉到僕人家裏過夜，洗你們的腳，清早起來再上路。」他們說：「不！我們要在廣場上過夜。」
GEN|19|3|羅得 懇切地請他們，他們就轉向他，進到他屋裏。 羅得 為他們預備宴席，烤無酵餅，他們就吃了。
GEN|19|4|他們還沒有躺下， 所多瑪城 的人，連老帶少所有的人，個個都來圍住那屋子。
GEN|19|5|他們呼叫 羅得 ，對他說：「今天晚上到你這裏來的人在哪裏？把他們帶出來，讓我們親近他們。」
GEN|19|6|羅得 出了門，把身後的門關上，到眾人那裏，
GEN|19|7|說：「我的弟兄們，請你們不要做這惡事。
GEN|19|8|看哪，我有兩個女兒，還沒有親近過男人，讓我領她們出來給你們，就照你們看為好的對待她們吧！只是這兩個人既然到我舍下，請不要向他們做這事。」
GEN|19|9|眾人說：「站到一邊去吧！」又說：「這個人來寄居，還想扮審判官呢！現在我們要害你比害他們更厲害。」眾人就往前衝向 羅得 ，要攻破大門。
GEN|19|10|那兩個人伸出手來，把 羅得 拉進屋子他們那裏，就關上門。
GEN|19|11|他們擊打門外的人，無論老少，都眼睛迷糊，找門找得很煩躁。
GEN|19|12|那兩個人對 羅得 說：「你這裏還有甚麼人嗎？無論是女婿，是兒女，這城中所有屬你的人，你都要把他們從這地方帶出去。
GEN|19|13|我們要毀滅這地方，因為控告城內百姓的聲音在耶和華面前非常大，耶和華派我們來毀滅這城。」
GEN|19|14|羅得 出去，告訴娶了 他女兒的女婿們說：「起來，離開這地方，因為耶和華要毀滅這城。」他的女婿們卻以為他說的是笑話。
GEN|19|15|天亮了，天使催逼 羅得 說：「起來！帶著你的妻子和你這裏的兩個女兒出去，免得你因這城的罪孽同被剿滅。」
GEN|19|16|但 羅得 遲延不走。二人因為耶和華憐憫 羅得 ，就拉著他的手和他妻子的手，以及他兩個女兒的手，把他們領出來，安置在城外；
GEN|19|17|領他們出來以後，就說：「逃命吧！不可回頭看，也不可在平原站住。要往山上逃跑，免得你被剿滅。」
GEN|19|18|羅得 對他們說：「我主啊，不要這樣！
GEN|19|19|看哪，你僕人已經在你眼前蒙恩，你又向我大施慈愛，救我的性命。但是我不能逃到山上去，恐怕這災禍追上我，我就死了。
GEN|19|20|看哪，這城又近又小，比較容易逃到那裏。這不是一座小城嗎？求你容我逃到那裏，使我的性命可以存活。」
GEN|19|21|天使對他說：「看哪，這事我也應允你，不傾覆你所說的這城。
GEN|19|22|你要趕快逃到那城，因為你還沒有到那裏，我不能做甚麼。」因此那城名叫 瑣珥 。
GEN|19|23|羅得 到了 瑣珥 ，太陽已經升出地面。
GEN|19|24|當時，耶和華把硫磺與火，從天上耶和華那裏降與 所多瑪 和 蛾摩拉 ，
GEN|19|25|把那些城和全平原，城裏所有的居民和土地上生長的，都毀滅了。
GEN|19|26|羅得 的妻子在他後邊回頭一看，就變成了一根鹽柱。
GEN|19|27|亞伯拉罕 清早起來，到了他先前站在耶和華面前的地方，
GEN|19|28|面向 所多瑪 和 蛾摩拉 ，以及平原全地觀望。他觀看，看哪，那地有濃煙上騰，好像燒窯的濃煙。
GEN|19|29|當上帝毀滅平原諸城的時候，他記念 亞伯拉罕 ；在傾覆 羅得 所住之城的時候，就把 羅得 從傾覆中帶出來。
GEN|19|30|羅得 因為怕住在 瑣珥 ，就同他兩個女兒從 瑣珥 上去，住在山上。他和兩個女兒住在一個洞裏。
GEN|19|31|大女兒對小女兒說：「我們的父親老了，這地又沒有男人可以照世上的禮俗來與我們結合。
GEN|19|32|來！我們叫父親喝酒，然後與他同寢。這樣，我們可以從我們的父親存留後裔。」
GEN|19|33|於是，那晚她們叫父親喝酒，大女兒就進去和她父親同寢；她幾時躺下，幾時起來，父親都不知道。
GEN|19|34|第二天，大女兒對小女兒說：「看哪，我昨夜與父親同寢。今晚我們再叫他喝酒，你進去與他同寢。這樣，我們可以從父親存留後裔。」
GEN|19|35|於是，那晚她們又叫父親喝酒，小女兒起來與她父親同寢；她幾時躺下，幾時起來，父親都不知道。
GEN|19|36|這樣， 羅得 的兩個女兒都從她們的父親懷了孕。
GEN|19|37|大女兒生了兒子，給他起名叫 摩押 ，就是現今 摩押 人的始祖。
GEN|19|38|小女兒也生了兒子，給他起名叫 便‧亞米 ，就是現今 亞捫 人的始祖。
GEN|20|1|亞伯拉罕 從那裏往 尼革夫 遷移，寄居在 加低斯 和 書珥 之間的 基拉耳 。
GEN|20|2|亞伯拉罕 稱他的妻子 撒拉 為妹妹。 基拉耳 王 亞比米勒 派人把 撒拉 帶走。
GEN|20|3|夜間，上帝在夢中來到 亞比米勒 那裏，對他說：「看哪，你要死了，因為你帶來的女人，她是有丈夫的女子！」
GEN|20|4|亞比米勒 還未親近 撒拉 ；他說：「主啊，連公義的國，你也要毀滅嗎？
GEN|20|5|那人豈不是自己對我說『她是我妹妹』嗎？連這女人自己也說：『他是我哥哥。』我做這事是心正手潔的。」
GEN|20|6|上帝在夢中對他說：「我也知道你做這事是心中正直的；是我攔阻了你，免得你得罪我。所以我不讓你侵犯她。
GEN|20|7|現在你當把這人的妻子歸還給他；因為他是先知，他要為你禱告，使你存活。你若不歸還，你當知道，你和你所有的人都必定死。」
GEN|20|8|亞比米勒 清早起來，叫了他的眾臣僕來，把這一切事說給他們聽，他們就很害怕。
GEN|20|9|亞比米勒 召了 亞伯拉罕 來，對他說：「你怎麼向我這樣做呢？我甚麼事得罪你，你竟使我和我的國陷在大罪中呢？你對我做了不該做的事了！」
GEN|20|10|亞比米勒 對 亞伯拉罕 說：「你看見甚麼才做這事呢？」
GEN|20|11|亞伯拉罕 說：「我以為這地方的人根本不敬畏上帝，必為我妻子的緣故殺我。
GEN|20|12|況且她也真是我的妹妹；她與我是同父異母的，後來作了我的妻子。
GEN|20|13|當上帝叫我離開父家、飄流在外的時候，我對她說：我們無論走到甚麼地方，你要對人說：『他是我哥哥』，這就是你以慈愛待我了。」
GEN|20|14|亞比米勒 把牛、羊、奴僕、婢女送給 亞伯拉罕 ，也把他的妻子 撒拉 歸還給他。
GEN|20|15|亞比米勒 說：「看哪，我的地都在你面前，你看為好的地方就居住吧。」
GEN|20|16|他對 撒拉 說：「看哪，我給你哥哥一千銀子。看哪，這要在你全家人面前遮羞 ，向眾人證實你是清白的。」
GEN|20|17|亞伯拉罕 向上帝禱告，上帝就醫好 亞比米勒 和他的妻子，以及他的使女們，他們就能生育。
GEN|20|18|因耶和華為 亞伯拉罕 的妻子 撒拉 的緣故，已經使 亞比米勒 家中的婦人不能懷孕。
GEN|21|1|耶和華照著他所說的眷顧 撒拉 ，耶和華實現了他對 撒拉 的應許。
GEN|21|2|亞伯拉罕 年老，到上帝對他說的那所定的時候， 撒拉 懷了孕，給他生了一個兒子。
GEN|21|3|亞伯拉罕 給 撒拉 所生的兒子起名叫 以撒 。
GEN|21|4|以撒 出生後第八日， 亞伯拉罕 遵照上帝所吩咐的，為 以撒 行割禮。
GEN|21|5|他兒子 以撒 出生的時候， 亞伯拉罕 年一百歲。
GEN|21|6|撒拉 說：「上帝使我歡笑，凡聽見的人必與我一同歡笑」，
GEN|21|7|又說：「誰能預先對 亞伯拉罕 說， 撒拉 要乳養孩子呢？因為在他年老的時候，我為他生了一個兒子。」
GEN|21|8|孩子漸漸長大，就斷了奶。 以撒 斷奶的那一天， 亞伯拉罕 擺設豐盛的宴席。
GEN|21|9|那時， 撒拉 看見 埃及 人 夏甲 為 亞伯拉罕 所生的兒子戲笑，
GEN|21|10|就對 亞伯拉罕 說：「你把這使女和她兒子趕出去！因為這使女的兒子不可與我的兒子 以撒 一同承受產業。」
GEN|21|11|亞伯拉罕 為這事非常憂愁，因為關乎他的兒子。
GEN|21|12|上帝對 亞伯拉罕 說：「你不必為這孩子和你的使女憂愁。 撒拉 對你說的話，你都要聽從；因為從 以撒 生的，才要稱為你的後裔。
GEN|21|13|至於使女的兒子，我也必使他成為一國，因為他是你的後裔。」
GEN|21|14|亞伯拉罕 清早起來，拿餅和一皮袋水，給了 夏甲 ，搭在她肩上，把她和孩子一起送走。 夏甲 就走了，但她卻在 別是巴 的曠野流浪。
GEN|21|15|皮袋的水用完了， 夏甲 就把孩子放在一棵小樹下，
GEN|21|16|自己走開約有一箭之遠，相對而坐，說：「我不忍心看見孩子死」。她就坐在對面，放聲大哭。
GEN|21|17|上帝聽見孩子的聲音，上帝的使者就從天上呼叫 夏甲 說：「 夏甲 ，你為何這樣呢？不要害怕，上帝已經聽見孩子在那裏的聲音了。
GEN|21|18|起來！把孩子扶起來，用你的手握住他，因我必使他成為大國。」
GEN|21|19|上帝開了 夏甲 的眼睛，她就看見一口水井。她就去，把皮袋裝滿了水，給孩子喝。
GEN|21|20|上帝與這孩子同在，他就漸漸長大，住在曠野，成了一個弓箭手。
GEN|21|21|他住在 巴蘭 的曠野；他母親從 埃及 地為他娶了一個妻子。
GEN|21|22|那時候， 亞比米勒 和他的將軍 非各 對 亞伯拉罕 說：「凡你所做的事，上帝都與你同在。
GEN|21|23|我願你如今在這裏指著上帝對我起誓，不要虧待我和我的兒子，以及我的子孫。我怎樣忠誠待你，你也要照樣忠誠待我和你所寄居的這地。」
GEN|21|24|亞伯拉罕 說：「我願意起誓。」
GEN|21|25|先前， 亞比米勒 的僕人霸佔了一口水井， 亞伯拉罕 為這事責備 亞比米勒 。
GEN|21|26|亞比米勒 說：「我不知道誰做了這事，你也沒有告訴我，我到今日才聽到。」
GEN|21|27|亞伯拉罕 把羊和牛給了 亞比米勒 ，二人就彼此立約。
GEN|21|28|亞伯拉罕 把七隻小母羊另放在一處。
GEN|21|29|亞比米勒 對 亞伯拉罕 說：「你把這七隻小母羊另放一處是甚麼意思呢？」
GEN|21|30|他說：「你要從我手裏接受這七隻小母羊，作我挖了這口井的證據。」
GEN|21|31|所以他給那地方起名叫 別是巴 ，因為他們二人在那裏起了誓。
GEN|21|32|他們在 別是巴 立了約， 亞比米勒 就和他的將軍 非各 起身回 非利士 人的地去了。
GEN|21|33|亞伯拉罕 就在 別是巴 種了一棵柳樹，在那裏求告耶和華—永恆上帝的名。
GEN|21|34|亞伯拉罕 在 非利士 人的地寄居了許多日子。
GEN|22|1|這些事以後，上帝考驗 亞伯拉罕 ，對他說：「 亞伯拉罕 ！」他說：「我在這裏。」
GEN|22|2|上帝說：「你要帶你的兒子，就是你所愛的獨子 以撒 ，往 摩利亞 地去，在我指示你的一座山上，把他獻為燔祭。」
GEN|22|3|亞伯拉罕 清早起來，預備了驢，帶著跟他一起的兩個僕人和他兒子 以撒 ，劈好了燔祭的柴，就起身往上帝指示他的地方去了。
GEN|22|4|到了第三日， 亞伯拉罕 舉目遙望那地方。
GEN|22|5|亞伯拉罕 對他的僕人說：「你們和驢留在這裏，我和孩子要去那裏敬拜，然後回到你們這裏來。」
GEN|22|6|亞伯拉罕 把燔祭的柴放在他兒子 以撒 身上，自己手裏拿著火與刀；於是二人同行。
GEN|22|7|以撒 對他父親 亞伯拉罕 說：「我父啊！」 亞伯拉罕 說：「我兒，我在這裏。」 以撒 說：「看哪，火與柴都有了，但燔祭的羔羊在哪裏呢？」
GEN|22|8|亞伯拉罕 說：「我兒，上帝必自己預備燔祭的羔羊。」於是二人同行。
GEN|22|9|他們到了上帝指示他的地方， 亞伯拉罕 在那裏築壇，把柴擺好，綁了他兒子 以撒 ，放在壇的柴上。
GEN|22|10|亞伯拉罕 就伸手拿刀，要殺他的兒子。
GEN|22|11|耶和華的使者從天上呼喚他說：「 亞伯拉罕 ！ 亞伯拉罕 ！」他說：「我在這裏。」
GEN|22|12|天使說：「不可在這孩子身上下手！一點也不可傷害他！現在我知道你是敬畏上帝的人了，因為你沒有把你的兒子，就是你的獨子，留下不給我。」
GEN|22|13|亞伯拉罕 舉目觀看，看哪，一隻公綿羊兩角纏在灌木叢中。 亞伯拉罕 就去牽了那隻公綿羊，獻為燔祭，代替他的兒子。
GEN|22|14|亞伯拉罕 給那地方起名叫「耶和華以勒」 。直到今日人還說：「在耶和華的山上必有預備。」
GEN|22|15|耶和華的使者第二次從天上呼喚 亞伯拉罕 ，
GEN|22|16|說：「耶和華說：『你既行了這事，沒有留下你的兒子，就是你的獨子，我指著自己起誓：
GEN|22|17|我必多多賜福給你，我必使你的後裔大大增多，如同天上的星、海邊的沙。你的後裔必得仇敵的城門，
GEN|22|18|並且地上的萬國都必因你的後裔得福，因為你聽從了我的話。』」
GEN|22|19|於是 亞伯拉罕 回到他僕人那裏。他們一同起身，往 別是巴 去， 亞伯拉罕 就住在 別是巴 。
GEN|22|20|這些事以後，有人告訴 亞伯拉罕 說：「看哪， 密迦 也為你兄弟 拿鶴 生了幾個兒子：
GEN|22|21|長子 烏斯 、他的兄弟 布斯 、 亞蘭 的父親 基摩利 、
GEN|22|22|基薛 、 哈瑣 、 必達 、 益拉 和 彼土利 。」
GEN|22|23|彼土利 生 利百加 。這八個人都是 密迦 為 亞伯拉罕 的兄弟 拿鶴 生的。
GEN|22|24|拿鶴 的妾名叫 流瑪 ，她也生了 提八 、 迦含 、 他轄 和 瑪迦 。
GEN|23|1|撒拉 享壽一百二十七歲，這是 撒拉 一生的歲數 。
GEN|23|2|撒拉 死在 迦南 地的 基列‧亞巴 ，就是 希伯崙 。 亞伯拉罕 來哀悼 撒拉 ，為她哭泣。
GEN|23|3|然後， 亞伯拉罕 起來，離開死人面前，對 赫 人說：
GEN|23|4|「我在你們中間是外人，是寄居的。請給我你們那裏的一塊墳地，我好埋葬我的亡妻，使她不在我的面前。」
GEN|23|5|赫 人回答 亞伯拉罕 說：
GEN|23|6|「我主請聽。你在我們中間是一位尊貴的王子，只管在我們最好的墳地裏埋葬你的死人；我們沒有一人會拒絕你在他的墳地裏埋葬你的死人。」
GEN|23|7|於是， 亞伯拉罕 起來，向當地的百姓 赫 人下拜，
GEN|23|8|對他們說：「你們若願意讓我埋葬我的亡妻，使她不在我面前，就請聽我，為我求 瑣轄 的兒子 以弗崙 ，
GEN|23|9|把他田地盡頭的 麥比拉洞 賣給我。他可以按照足價賣給我，作為我在你們中間的墳地。」
GEN|23|10|那時， 以弗崙 正坐在 赫 人中間。 赫 人 以弗崙 就回答 亞伯拉罕 ，說給所有出入城門的 赫 人聽：
GEN|23|11|「不，我主請聽。我要把這塊田送給你，連田間的洞也送給你，在我同族的人眼前都給你，讓你埋葬你的死人。」
GEN|23|12|亞伯拉罕 就在當地的百姓面前下拜，
GEN|23|13|對 以弗崙 說，也給當地百姓聽：「你若應允，請你聽我。我要把田的價錢給你，請你收下，我就在那裏埋葬我的死人。」
GEN|23|14|以弗崙 回答 亞伯拉罕 說：
GEN|23|15|「我主請聽。四百舍客勒銀子的地，在你我中間算甚麼呢？只管埋葬你的死人吧！」
GEN|23|16|亞伯拉罕 聽從了 以弗崙 。 亞伯拉罕 就照著他說給 赫 人聽的，把買賣通用的銀子，秤了四百舍客勒銀子給 以弗崙 。
GEN|23|17|於是， 以弗崙 把那塊位於 幔利 對面的 麥比拉 田，和其中的洞，以及田間周圍的樹木都成交了，
GEN|23|18|在所有出入城門的 赫 人眼前，賣給 亞伯拉罕 作為他的產業。
GEN|23|19|後來， 亞伯拉罕 把他妻子 撒拉 安葬在 迦南 地 幔利 對面的 麥比拉 田間的洞裏， 幔利 就是 希伯崙 。
GEN|23|20|從此，那塊田和田間的洞就從 赫 人移交給 亞伯拉罕 作墳地的產業。
GEN|24|1|亞伯拉罕 年紀老邁，耶和華在一切事上都賜福給他。
GEN|24|2|亞伯拉罕 對他家中管理他一切產業最老的僕人說：「把你的手放在我大腿底下。
GEN|24|3|我要叫你指著耶和華—天和地的上帝起誓，不要為我兒子娶我所居住的 迦南 地的女子為妻。
GEN|24|4|你要往我的本地本族去，為我的兒子 以撒 娶妻。」
GEN|24|5|僕人對他說：「如果那女子不肯跟我來到這地，我必須把你的兒子帶回到你出來的地方嗎？」
GEN|24|6|亞伯拉罕 對他說：「你要謹慎，不可帶我兒子回那裏去。
GEN|24|7|耶和華—天上的上帝曾帶領我離開父家和本族的地，對我說話，向我起誓說：『我要將這地賜給你的後裔。』他要差遣使者在你面前，你就可以從那裏為我兒子娶妻。
GEN|24|8|倘若那女子不肯跟你來，我叫你起的誓就與你無關了，只是你不可帶我的兒子回到那裏去。」
GEN|24|9|僕人就把手放在他主人 亞伯拉罕 的大腿底下，為這事向他起誓。
GEN|24|10|那僕人從他主人的駱駝中取了十匹駱駝，他手中也帶著他主人各樣的貴重物品離開 ，起身往 美索不達米亞 去，到了 拿鶴 的城。
GEN|24|11|傍晚時，眾女子出來打水，他就讓駱駝跪在城外的水井旁。
GEN|24|12|他說：「耶和華—我主人 亞伯拉罕 的上帝啊，求你施恩給我的主人 亞伯拉罕 ，讓我今日就遇見吧！
GEN|24|13|看哪，我站在井旁，城內居民的女子們正出來打水。
GEN|24|14|我向哪一個少女說：『請你放下水瓶來，給我水喝』，她若說：『請喝！我也給你的駱駝喝』，願她作你所選定給你僕人 以撒 的妻。這樣，我就知道你施恩給我的主人了。」
GEN|24|15|話還沒說完，看哪， 利百加 肩頭上扛著水瓶出來。 利百加 是 彼土利 所生的； 彼土利 是 亞伯拉罕 的兄弟 拿鶴 妻子 密迦 的兒子。
GEN|24|16|那少女容貌極其美麗，是未曾與人親近的童女。她下到井旁，打滿了瓶子的水，就上來。
GEN|24|17|僕人跑上前去迎著她，說：「請你讓我喝你瓶子裏的一點水。」
GEN|24|18|少女說：「我主請喝！」就急忙拿下瓶子托在手上，給他喝水。
GEN|24|19|那少女給他喝足了，又說：「我也為你的駱駝打水，直到駱駝喝足了。」
GEN|24|20|她就急忙把瓶子裏的水倒在槽裏，又跑到井旁打水，為所有的駱駝打了水。
GEN|24|21|那人定睛看著少女，一句話也不說，要知道耶和華是否使他的道路亨通。
GEN|24|22|駱駝喝足了，那人就拿出一個比加 重的金環，一對十舍客勒重的金手鐲，
GEN|24|23|說：「請告訴我，你是誰的女兒？你父親家裏有沒有地方可以讓我們過夜？」
GEN|24|24|少女說：「我是 密迦 為 拿鶴 生的兒子 彼土利 的女兒。」
GEN|24|25|又說：「我們家裏有充足的乾草和飼料，也有住宿的地方。」
GEN|24|26|那人就低頭向耶和華敬拜，
GEN|24|27|說：「耶和華—我主人 亞伯拉罕 的上帝是應當稱頌的，因他不斷以慈愛信實待我主人。至於我，耶和華一路引領我，直到我主人的兄弟家裏。」
GEN|24|28|那少女跑去，把這些話告訴她母親家裏的人。
GEN|24|29|利百加 有一個哥哥，名叫 拉班 ， 拉班 就跑到外面井旁那人那裏。
GEN|24|30|當他看見金環和戴在他妹妹手上的金鐲，又聽見他妹妹 利百加 說的話：「那人如此對我說」，他就來到那人面前，看哪，他還站在井旁的駱駝旁邊，
GEN|24|31|就對他說：「你這蒙耶和華賜福的人，請進來吧！為甚麼站在外面？我已經收拾了房屋，也為駱駝預備了地方。」
GEN|24|32|那人就進了 拉班 的家。 拉班 卸了駱駝，用飼料餵牠們，拿水給那人和隨從他的人洗腳，
GEN|24|33|把食物擺在他面前，請他吃。他卻說：「我不吃，等我把我的事情說完了再吃。」 拉班 說：「請說。」
GEN|24|34|他說：「我是 亞伯拉罕 的僕人。
GEN|24|35|耶和華大大地賜福給我主人，使他發達，賜給他羊群、牛群、金銀、奴僕、婢女、駱駝和驢。
GEN|24|36|我主人的妻子 撒拉 年老的時候為我主人生了一個兒子；我主人把他一切所有的都給了他。
GEN|24|37|我主人叫我起誓說：『不要為我兒子娶我所居住的 迦南 地的女子為妻。
GEN|24|38|你要往我父家、我本族那裏去，為我的兒子娶妻。』
GEN|24|39|我對我主人說：『恐怕那女子不肯跟我來。』
GEN|24|40|他就說：『我所事奉的耶和華必要差遣他的使者與你同去，使你的道路亨通，你就可以在我父家、我本族那裏，為我的兒子娶妻。
GEN|24|41|只要你到了我本族那裏，我叫你起的誓就與你無關。他們若不把女子交給你，我叫你起的誓也與你無關。』
GEN|24|42|「我今日到了井旁，就說：『耶和華—我主人 亞伯拉罕 的上帝啊，願你使我所行的道路亨通。
GEN|24|43|看哪，我站在井旁，對哪一個出來打水的女子說：請你讓我喝你瓶子裏的一點水，
GEN|24|44|她若說：你只管喝，我也為你的駱駝打水；願那女子作耶和華給我主人兒子所選定的妻子。』
GEN|24|45|「我心裏的話還沒有說完，看哪， 利百加 肩頭上扛著水瓶出來，下到井旁打水。我對她說：『請你給我水喝。』
GEN|24|46|她就急忙從肩頭上拿下瓶子來，說：『請喝！我也給你的駱駝喝。』我就喝了；她也給我的駱駝喝了。
GEN|24|47|我問她說：『你是誰的女兒？』她說：『我是 彼土利 的女兒， 彼土利 是 密迦 和 拿鶴 生的兒子。』我就把環子戴在她鼻子上，把鐲子戴在她雙手上。
GEN|24|48|然後我低頭向耶和華敬拜，稱頌耶和華—我主人 亞伯拉罕 的上帝，因為他引導我走合適的道路，使我得著我主人兄弟的孫女，給我主人的兒子為妻。
GEN|24|49|現在你們若願以慈愛誠信待我主人，就告訴我；若不然，也告訴我，使我可以或向左，或向右。」
GEN|24|50|拉班 和 彼土利 回答說：「這事既然出於耶和華，我們不能向你說好說歹。
GEN|24|51|看哪， 利百加 就在你面前，可以將她帶去，遵照耶和華所說的，給你主人的兒子為妻。」
GEN|24|52|亞伯拉罕 的僕人聽見他們這些話，就向耶和華俯伏在地。
GEN|24|53|僕人拿出金器、銀器和衣服送給 利百加 ，又將貴重的物品送給她哥哥和她母親。
GEN|24|54|然後，僕人和隨從的人才吃喝，並且住了一夜。早晨起來，僕人說：「請讓我回我主人那裏去吧。」
GEN|24|55|利百加 的哥哥和母親說：「讓她同我們再住幾天，也許十天，然後她可以去。」
GEN|24|56|僕人對他們說：「耶和華既然使我道路亨通，你們就不要耽誤我，請讓我走，回我主人那裏去吧！」
GEN|24|57|他們說：「我們把她叫來問問她 。」
GEN|24|58|他們就叫了 利百加 來，對她說：「你和這人同去嗎？」她說：「我去。」
GEN|24|59|於是他們送他們的妹妹 利百加 和她的奶媽，同 亞伯拉罕 的僕人，以及隨從他的人走了。
GEN|24|60|他們就為 利百加 祝福，對她說： 「我們的妹妹啊， 願你作千萬人的母親！ 願你的後裔得著仇敵的城門！」
GEN|24|61|利百加 和她的女僕們起來，騎上駱駝，跟著那人去。僕人就帶著 利百加 走了。
GEN|24|62|那時， 以撒 住在 尼革夫 。他剛從 庇耳‧拉海‧萊 回來。
GEN|24|63|傍晚時， 以撒 出來，到田間默想。他舉目一看，看哪，來了一隊駱駝。
GEN|24|64|利百加 舉目看見 以撒 ，就急忙下了駱駝，
GEN|24|65|對那僕人說：「這從田間走來迎接我們的人是誰？」僕人說：「他是我的主人。」 利百加 就拿面紗蓋住自己。
GEN|24|66|僕人把他所做的一切事都告訴 以撒 。
GEN|24|67|以撒 就領 利百加 進了母親 撒拉 的帳棚，娶了她為妻，並且愛她。 以撒 自從母親離世以後，這才得了安慰。
GEN|25|1|亞伯拉罕 再娶了一個妻子，名叫 基土拉 。
GEN|25|2|她為他生了 心蘭 、 約珊 、 米但 、 米甸 、 伊施巴 和 書亞 。
GEN|25|3|約珊 生了 示巴 和 底但 。 底但 的子孫是 亞書利 族、 利都是 族和 利烏米 族。
GEN|25|4|米甸 的兒子是 以法 、 以弗 、 哈諾 、 亞比大 和 以勒大 。這些都是 基土拉 的子孫。
GEN|25|5|亞伯拉罕 把他一切所有的都給了 以撒 。
GEN|25|6|至於 亞伯拉罕 妾的兒子， 亞伯拉罕 趁著自己還活著的時候把財物分給他們，打發他們離開他的兒子 以撒 ，往東方去，直到東方之地。
GEN|25|7|這是 亞伯拉罕 一生的年日，他活了一百七十五年。
GEN|25|8|亞伯拉罕 壽高年邁，安享天年，息勞而終，歸到他祖先 那裏。
GEN|25|9|他兩個兒子 以撒 、 以實瑪利 把他安葬在 麥比拉 洞裏。這洞在 幔利 的對面、 赫 人 瑣轄 的兒子 以弗崙 的田中，
GEN|25|10|就是 亞伯拉罕 向 赫 人買的那塊田。 亞伯拉罕 和他妻子 撒拉 都葬在那裏。
GEN|25|11|亞伯拉罕 死了以後，上帝賜福給他的兒子 以撒 。 以撒 住在 庇耳‧拉海‧萊 附近。
GEN|25|12|這是 撒拉 的婢女、 埃及 人 夏甲 為 亞伯拉罕 生的兒子 以實瑪利 的後代。
GEN|25|13|以實瑪利 兒子們的名字，按著他們後代的名字如下： 以實瑪利 的長子 尼拜約 ，又有 基達 、 亞德別 、 米比衫 、
GEN|25|14|米施瑪 、 度瑪 、 瑪撒 、
GEN|25|15|哈大 、 提瑪 、 伊突 、 拿非施 ，和 基底瑪 。
GEN|25|16|這些都是 以實瑪利 的兒子們。他們的村莊和營寨按著他們命名；他們作了十二族的族長。
GEN|25|17|以實瑪利 一生的歲數是一百三十七歲，斷氣而死，歸到他祖先那裏。
GEN|25|18|他的子孫住在 哈腓拉 ，直到 埃及 東邊的 書珥 ，向著 亞述 ，在他眾弟兄的對面安頓下來 。
GEN|25|19|這是 亞伯拉罕 的兒子 以撒 的後代。 亞伯拉罕 生 以撒 。
GEN|25|20|以撒 四十歲時娶 利百加 為妻。 利百加 是 巴旦‧亞蘭 地的 亞蘭 人 彼土利 的女兒，是 亞蘭 人 拉班 的妹妹。
GEN|25|21|以撒 因他妻子不生育，就為她祈求耶和華。耶和華應允他的祈求，他的妻子 利百加 就懷了孕。
GEN|25|22|胎兒們在她腹中彼此相爭，她就說：「若是如此，我為甚麼會這樣呢 ？」她就去求問耶和華。
GEN|25|23|耶和華對她說： 兩國在你腹中； 兩族要從你身上分立。 這族必強於那族； 將來大的要服侍小的。
GEN|25|24|到了生產的日期，看哪，腹中是對雙胞胎。
GEN|25|25|先出生的身體帶紅，渾身有毛，好像皮衣；他們就給他起名叫 以掃 。
GEN|25|26|隨後， 以掃 的弟弟也出生，他的手抓住 以掃 的腳跟，因此給他起名叫 雅各 。兩個兒子出生時， 以撒 六十歲。
GEN|25|27|兩個孩子漸漸長大， 以掃 善於打獵，常在田野； 雅各 為人安靜，常住在帳棚裏。
GEN|25|28|以撒 愛 以掃 ，因為常吃他的野味； 利百加 卻愛 雅各 。
GEN|25|29|有一天， 雅各 熬了湯， 以掃 從田野回來，疲憊不堪。
GEN|25|30|以掃 對 雅各 說：「我累死了，請你讓我吃這紅的，這紅的湯吧！」因此 以掃 又叫 以東 。
GEN|25|31|雅各 說：「你今日把長子的名分賣給我吧。」
GEN|25|32|以掃 說：「看哪，我快要死了，這長子的名分對我有甚麼用呢？」
GEN|25|33|雅各 說：「你今日對我起誓吧。」 以掃 就向他起誓，把長子的名分賣給了 雅各 。
GEN|25|34|於是 雅各 把餅和豆湯給了 以掃 ， 以掃 吃喝以後，起來走了。這樣， 以掃 輕看他長子的名分。
GEN|26|1|那地有了饑荒，不是 亞伯拉罕 的時候曾有過的那次饑荒， 以撒 就到 基拉耳 ， 非利士 人的王 亞比米勒 那裏去。
GEN|26|2|耶和華向 以撒 顯現，說：「你不要下 埃及 去，要住在我所指示你的地。
GEN|26|3|你要寄居在這地，我必與你同在，賜福給你，因為我要將這一切的地都賜給你和你的後裔。我必堅定我向你父親 亞伯拉罕 所起的誓。
GEN|26|4|我要使你的後裔增多，好像天上的星，又要將這一切的地賜給你的後裔，並且地上的萬國都必因你的後裔得福，
GEN|26|5|因為 亞伯拉罕 聽從我的話，遵守我的吩咐、誡令、律例和教導。」
GEN|26|6|於是， 以撒 住在 基拉耳 。
GEN|26|7|那地方的人問起他的妻子，他就說：「她是我的妹妹。」原來他害怕說「我的妻子」。他想：「或許這地方的人會因 利百加 殺我，因為她容貌美麗。」
GEN|26|8|他在那裏住了一段很長的日子。有一天， 非利士 人的王 亞比米勒 從窗戶往外觀看，看哪， 以撒 在撫愛他的妻子 利百加 。
GEN|26|9|亞比米勒 召 以撒 來，說：「看哪，她實在是你的妻子，你怎麼說『她是我的妹妹』呢？」 以撒 對他說：「因為我想，恐怕我會因她而死。」
GEN|26|10|亞比米勒 說：「你向我們做的是甚麼事呢？百姓中有一個人幾乎要和你的妻子同寢，你就把我們陷在罪中了。」
GEN|26|11|於是 亞比米勒 命令眾百姓說：「凡侵犯這個人，或他妻子的，必要把他處死。」
GEN|26|12|以撒 在那地耕種，那一年有百倍的收成。耶和華賜福給他，
GEN|26|13|他就發達，日漸昌盛，成了大富翁。
GEN|26|14|他有羊群牛群，又有許多僕人， 非利士 人就嫉妒他。
GEN|26|15|他父親 亞伯拉罕 在世的時候，他父親的僕人所挖的井， 非利士 人全都塞住，填滿了土。
GEN|26|16|亞比米勒 對 以撒 說：「你離開我們去吧，因為你比我們強盛得多。」
GEN|26|17|以撒 就離開那裏，在 基拉耳谷 支搭帳棚，住在那裏。
GEN|26|18|他父親 亞伯拉罕 在世的時候所挖的水井，在 亞伯拉罕 死後，都被 非利士 人塞住了， 以撒 就重新把井挖出來，仍照他父親所取的名為它們命名。
GEN|26|19|以撒 的僕人在谷中挖井，就在那裏得了一口活水井。
GEN|26|20|基拉耳 的牧人與 以撒 的牧人相爭，說：「這水是我們的。」 以撒 就給那井起名叫 埃色 ，因為他們和他相爭。
GEN|26|21|以撒 的僕人又挖了一口井，他們又為這井相爭， 以撒 就給這井起名叫 西提拿 。
GEN|26|22|以撒 離開那裏，又挖了一口井，他們不再為這井相爭了，他就給那井起名叫 利河伯 。他說：「耶和華現在給我們寬闊之地，我們必在這地興旺。」
GEN|26|23|以撒 從那裏上 別是巴 去。
GEN|26|24|當夜耶和華向他顯現，說：「我是你父親 亞伯拉罕 的上帝。不要懼怕，因為我與你同在，要賜福給你，也要為我僕人 亞伯拉罕 的緣故，使你的後裔增多。」
GEN|26|25|以撒 就在那裏築了一座壇，求告耶和華的名，並且在那裏支搭帳棚；他的僕人就在那裏挖了一口井。
GEN|26|26|亞比米勒 同他的顧問 亞戶撒 和他軍隊的元帥 非各 ，從 基拉耳 來到 以撒 那裏。
GEN|26|27|以撒 對他們說：「你們既然恨我，趕我離開你們，為甚麼又到我這裏來呢？」
GEN|26|28|他們說：「我們明明看見耶和華與你同在；因此就說，讓我們雙方彼此起誓，我們跟你立約，
GEN|26|29|使你不加害我們，正如我們未曾侵犯你，素來善待你，並且送你平平安安地走。你是蒙耶和華賜福的！」
GEN|26|30|以撒 為他們擺設宴席，他們就一起吃喝。
GEN|26|31|他們清早起來，彼此起誓。 以撒 送他們走，他們就平平安安地離開他去了。
GEN|26|32|那一天， 以撒 的僕人來，把挖井的消息告訴他，說：「我們得到水了。」
GEN|26|33|他就給那井起名叫 示巴 ，因此那城名叫 別是巴 ，直到今日。
GEN|26|34|以掃 四十歲的時候娶了 赫 人 比利 的女兒 猶滴 ，和 赫 人 以倫 的女兒 巴實抹 為妻。
GEN|26|35|她們使 以撒 和 利百加 心裏愁煩。
GEN|27|1|以撒 年老，眼睛昏花，不能看見，就叫他大兒子 以掃 來，對他說：「我兒。」 以掃 對他說：「我在這裏。」
GEN|27|2|他說：「看哪，我老了，不知道哪一天死。
GEN|27|3|現在拿你打獵的工具，就是箭囊和弓，到田野去為我打獵，
GEN|27|4|照我所愛的做成美味，拿來給我吃，好讓我在未死之前為你祝福。」
GEN|27|5|以撒 對他兒子 以掃 說話的時候， 利百加 聽見了。 以掃 往田野去打獵，要把獵物帶回來。
GEN|27|6|利百加 就對她兒子 雅各 說：「看哪，我聽見你父親對你哥哥 以掃 說：
GEN|27|7|『你去把獵物帶回來，做成美味給我吃，讓我在未死之前，在耶和華面前為你祝福。』
GEN|27|8|現在，我兒，你要聽我的話，照我所吩咐你的，
GEN|27|9|到羊群裏去，從那裏牽兩隻肥美的小山羊來給我，我就照你父親所愛的，把牠們做成美味給他。
GEN|27|10|然後，你拿到你父親那裏給他吃，好讓他在未死之前為你祝福。」
GEN|27|11|雅各 對他母親 利百加 說：「看哪，我哥哥 以掃 渾身都有毛，我身上卻是光滑的；
GEN|27|12|倘若父親摸著我，我在他眼中就是騙子了。這樣，我就自招詛咒，而不是祝福。」
GEN|27|13|他母親對他說：「我兒，你所受的詛咒臨到我身上吧！你只管聽我的話，去牽小山羊來給我。」
GEN|27|14|他就去牽來，交給他母親。他母親就照他父親所愛的，做成美味。
GEN|27|15|利百加 把大兒子 以掃 在家裏最好的衣服給她小兒子 雅各 穿，
GEN|27|16|又用小山羊的皮包在 雅各 的手上和頸項光滑的地方，
GEN|27|17|就把所做的美味和餅交在她兒子 雅各 的手裏。
GEN|27|18|雅各 來到他父親那裏，說：「我的父親！」他說：「我在這裏。我兒，你是誰？」
GEN|27|19|雅各 對他父親說：「我是你的長子 以掃 。我已照你吩咐我的做了。請起來坐著，吃我的野味，你好為我祝福。」
GEN|27|20|以撒 對他兒子說：「我兒，你怎麼這樣快就找到了呢？」他說：「因為這是耶和華—你的上帝使我遇見的。」
GEN|27|21|以撒 對 雅各 說：「我兒，靠近一點，讓我摸摸你，你真的是我的兒子 以掃 嗎？」
GEN|27|22|雅各 就靠近他父親 以撒 。 以撒 摸著他，說：「聲音是 雅各 的聲音，手卻是 以掃 的手。」
GEN|27|23|以撒 認不出他來，因為他手上有毛，像他哥哥 以掃 的手一樣。於是， 以撒 就為他祝福。
GEN|27|24|以撒 說：「你真的是我兒子 以掃 嗎？」他說：「我是。」
GEN|27|25|以撒 說：「拿給我，讓我吃我兒子的野味，我好為你祝福。」 雅各 拿給他，他就吃了，又拿酒給他，他也喝了。
GEN|27|26|他父親 以撒 對他說：「我兒，靠近一點來親我！」
GEN|27|27|他就近前親吻父親。他父親一聞他衣服上的香氣，就為他祝福，說： 「看，我兒的香氣 好像耶和華賜福之田地的香氣。
GEN|27|28|願上帝賜你天上的甘露， 地上的肥土， 和豐富的五穀新酒。
GEN|27|29|願萬民事奉你， 萬族向你下拜。 願你作你弟兄的主， 你母親的兒子向你下拜。 詛咒你的，願他受詛咒； 祝福你的，願他蒙祝福。」
GEN|27|30|以撒 為 雅各 祝福完畢， 雅各 才從他父親那裏出來，他哥哥 以掃 正打獵回來。
GEN|27|31|以掃 也做了美味，拿來給他父親，對他父親說：「父親，請起來，吃你兒子的野味，你好為我祝福。」
GEN|27|32|他父親 以撒 對他說：「你是誰？」他說：「我是你的兒子，你的長子 以掃 。」
GEN|27|33|以撒 就大大戰兢，說：「那麼，是誰打了獵物拿來給我呢？你未來之前我已經吃了，也為他祝福了，他將來就必蒙福。」
GEN|27|34|以掃 聽了他父親的話，就大聲痛哭，對他父親說：「我父啊，求你也為我祝福！」
GEN|27|35|以撒 說：「你弟弟已經用詭計來把你的福分奪去了。」
GEN|27|36|以掃 說：「他名叫 雅各 ，豈不是這樣嗎？他欺騙了我兩次：他先前奪了我長子的名分，看哪，他現在又奪了我的福分。」 以掃 又說：「你沒有留下給我的祝福嗎？」
GEN|27|37|以撒 回答 以掃 說：「看哪，我已立他作你的主，使他的弟兄都給他作僕人，並賜他五穀新酒可以養生。我兒，那麼，現在我還能為你做甚麼呢？」
GEN|27|38|以掃 對他父親說：「我父啊，你只有一個祝福嗎？我父啊，求你也為我祝福！」 以掃 就放聲而哭。
GEN|27|39|他父親 以撒 回答說： 「看哪，你所住的地方必缺乏肥沃的土地， 缺乏天上的甘露 。
GEN|27|40|你必倚靠刀劍度日， 又必服侍你的兄弟； 到你強盛的時候， 必從你頸項上掙開他的軛。
GEN|27|41|以掃 因他父親給 雅各 的祝福，就怨恨 雅各 ，心裏說：「為我父親居喪的時候近了，到那時候，我要殺我的弟弟 雅各 。」
GEN|27|42|有人把 利百加 大兒子 以掃 的話告訴 利百加 ，她就派人去，叫了她小兒子 雅各 來，對他說：「看哪，你哥哥 以掃 想要殺你來洩恨。
GEN|27|43|現在，我兒，聽我的話，起來，逃往 哈蘭 ，到我哥哥 拉班 那裏去，
GEN|27|44|同他住一段日子，直等到你哥哥的怒氣消了。
GEN|27|45|等到你哥哥向你消了怒氣，忘了你向他所做的事，我就派人去，把你從那裏帶回來。我何必在一天之內喪失你們二人呢？」
GEN|27|46|利百加 對 以撒 說：「我因這 赫 人的女子活得不耐煩了；倘若 雅各 也從本地女子中娶像這樣的 赫 人女子為妻，我為甚麼要活著呢？」
GEN|28|1|以撒 叫了 雅各 來，為他祝福，並吩咐他說：「你不要娶 迦南 的女子為妻。
GEN|28|2|你起身往 巴旦‧亞蘭 去，到你外祖父 彼土利 的家，從你舅父 拉班 的女兒中娶一位作你的妻子。
GEN|28|3|願全能的上帝賜福給你，使你生養眾多，成為許多民族，
GEN|28|4|將應許 亞伯拉罕 的福賜給你和你的後裔，使你承受你所寄居的地為業，就是上帝賜給 亞伯拉罕 的地。」
GEN|28|5|以撒 送 雅各 走了， 雅各 就往 巴旦‧亞蘭 去，到 亞蘭 人 彼土利 的兒子 拉班 那裏， 拉班 是 利百加 的哥哥， 利百加 是 雅各 和 以掃 的母親。
GEN|28|6|以掃 見 以撒 已經為 雅各 祝福，而且送他往 巴旦‧亞蘭 去，在那裏娶妻，並且見 以撒 祝福 雅各 的時候吩咐他說：「不要娶 迦南 的女子為妻」，
GEN|28|7|又見 雅各 聽從父母的話往 巴旦‧亞蘭 去了，
GEN|28|8|以掃 就看出他父親 以撒 看 迦南 女子不順眼。
GEN|28|9|於是他往 以實瑪利 那裏去，在兩個妻子之外， 又娶了 瑪哈拉 為妻，她是 亞伯拉罕 兒子 以實瑪利 的女兒，是 尼拜約 的妹妹。
GEN|28|10|雅各 離開 別是巴 ，往 哈蘭 去。
GEN|28|11|到了一個地方，因為已經日落，就在那裏過夜。他拾起那地方的一塊石頭枕在頭下，就躺在那地方。
GEN|28|12|他做夢，看哪，一個梯子立在地上，梯子的頂端直伸到天；看哪，上帝的使者在梯子上，上去下來。
GEN|28|13|看哪，耶和華站在梯子上面 ，說：「我是耶和華—你祖父 亞伯拉罕 的上帝， 以撒 的上帝。你現在躺臥之地，我要將它賜給你和你的後裔。
GEN|28|14|你的後裔必像地上的塵沙，必向東西南北開展；地上萬族必因你和你的後裔得福。
GEN|28|15|看哪，我必與你同在，無論你往哪裏去，我必保佑你，領你歸回這地。我總不離棄你，直到我實現了對你所說的話。」
GEN|28|16|雅各 睡醒了，說：「耶和華真的在這裏，我竟不知道！」
GEN|28|17|他就懼怕，說：「這地方何等可畏！這不是別的，是上帝的殿，是天的門。」
GEN|28|18|雅各 清早起來，拿起枕在頭下的石頭，立作柱子，澆油在上面。
GEN|28|19|他給那地方起名叫 伯特利 ；那地方原先名叫 路斯 。
GEN|28|20|雅各 許願說：「上帝若與我同在，在我所行的路上保佑我，給我食物吃，衣服穿，
GEN|28|21|使我平平安安回到我父親的家，我就必以耶和華為我的上帝。
GEN|28|22|我所立為柱子的這塊石頭必作上帝的殿；凡你所賜給我的，我必將十分之一獻給你。」
GEN|29|1|雅各 起行，到了東方人之地。
GEN|29|2|他觀看，看哪，田間有一口井，看哪，有三群羊臥在井旁；因為人都取那井裏的水給羊喝。井口上的那塊石頭很大。
GEN|29|3|羊群都在那裏聚集，人就把石頭移開井口，取水給羊喝，然後又把石頭放回井口原處。
GEN|29|4|雅各 對他們說：「弟兄們，你們從哪裏來？」他們說：「我們是從 哈蘭 來的。」
GEN|29|5|他對他們說：「你們認識 拿鶴 的孫子 拉班 嗎？」他們說：「我們認識。」
GEN|29|6|雅各 對他們說：「他平安嗎？」他們說：「平安。看哪，他女兒 拉結 和羊一起來了。」
GEN|29|7|雅各 說：「看哪，日正當中，不是牲畜聚集的時候。你們取水給羊喝，再去牧放吧！」
GEN|29|8|他們說：「我們不能這樣，必須等所有的羊群聚集，人把石頭移開井口，我們才可以取水給羊喝。」
GEN|29|9|雅各 正和他們說話的時候， 拉結 和她父親的羊來了，因為她是牧羊的。
GEN|29|10|雅各 看見他舅父 拉班 的女兒 拉結 和舅父 拉班 的羊群，就上前把石頭移開井口，取水給舅父 拉班 的羊喝。
GEN|29|11|雅各 親了 拉結 ，就放聲大哭。
GEN|29|12|雅各 告訴 拉結 ，自己是她父親的親戚 ，是 利百加 的兒子。 拉結 就跑去告訴她父親。
GEN|29|13|拉班 聽見外甥 雅各 的消息，就跑去迎接他，抱著他，親他，帶他到自己的家。 雅各 把這一切的事告訴 拉班 。
GEN|29|14|拉班 對他說：「你實在是我的骨肉。」 雅各 就和他同住了一個月。
GEN|29|15|拉班 對 雅各 說：「雖然你是我的親戚，怎麼可以讓你白白服事我呢？告訴我，你要甚麼作工資呢？」
GEN|29|16|拉班 有兩個女兒，大的名叫 利亞 ，小的名叫 拉結 。
GEN|29|17|利亞 的雙眼無神， 拉結 卻長得美貌秀麗。
GEN|29|18|雅各 愛 拉結 ，就說：「我願為你的小女兒 拉結 服事你七年。」
GEN|29|19|拉班 說：「我把她給你，勝過給別人，你與我同住吧！」
GEN|29|20|雅各 就為 拉結 服事了七年；他因為愛 拉結 ，就看這七年如同幾天。
GEN|29|21|雅各 對 拉班 說：「日期已經滿了，請把我的妻子給我，我好與她同房。」
GEN|29|22|拉班 就擺設宴席，請了當地所有的人。
GEN|29|23|到了晚上， 拉班 帶女兒 利亞 來送給 雅各 ， 雅各 就與她同房。
GEN|29|24|拉班 也把自己的婢女 悉帕 給女兒 利亞 作婢女。
GEN|29|25|到了早晨，看哪，她是 利亞 ， 雅各 對 拉班 說：「你向我做的是甚麼事呢？我服事你，不是為 拉結 嗎？你為甚麼欺騙我呢？」
GEN|29|26|拉班 說：「大女兒還沒有給人就先把小女兒給人，我們這地方沒有這樣的規矩。
GEN|29|27|你先為這個滿了七日，我們就把那個也給你，不過你要另外再服事我七年。」
GEN|29|28|雅各 就這樣做了。滿了 利亞 的七日， 拉班 就把女兒 拉結 給 雅各 為妻。
GEN|29|29|拉班 又把自己的婢女 辟拉 給女兒 拉結 作婢女。
GEN|29|30|雅各 也與 拉結 同房，並且愛 拉結 勝過愛 利亞 ，於是他又服事了 拉班 七年。
GEN|29|31|耶和華見 利亞 失寵 ，就使她生育， 拉結 卻不生育。
GEN|29|32|利亞 懷孕生子，給他起名叫 呂便 ，因為她說：「耶和華看見我的苦情，如今我的丈夫必愛我。」
GEN|29|33|她又懷孕生子，給他起名叫 西緬 ，說：「耶和華因為聽見我失寵，所以又賜給我這個兒子。」
GEN|29|34|她又懷孕生子，說：「我給丈夫生了三個兒子，現在，這次他必親近我了。」因此， 雅各 給他起名叫 利未 。
GEN|29|35|她又懷孕生子，說：「這次我要讚美耶和華。」因此給他起名叫 猶大 。於是她停了生育。
GEN|30|1|拉結 見自己不給 雅各 生孩子，就嫉妒她姊姊，對 雅各 說：「你給我孩子，不然，讓我死了吧。」
GEN|30|2|雅各 對 拉結 生氣，說：「是我代替上帝使你生不出孩子的嗎？」
GEN|30|3|拉結 說：「看哪，我的使女 辟拉 在這裏，你可以與她同房，使她生子歸在我膝下，我也可以藉著她得孩子 。」
GEN|30|4|拉結 就把她的婢女 辟拉 給丈夫為妾， 雅各 與她同房。
GEN|30|5|辟拉 懷孕，為 雅各 生了一個兒子。
GEN|30|6|拉結 給他起名叫 但 ，說：「上帝為我伸冤，也聽了我的聲音，賜給我一個兒子。」
GEN|30|7|拉結 的婢女 辟拉 又懷孕，為 雅各 生了第二個兒子。
GEN|30|8|拉結 給他起名叫 拿弗他利 ，說：「我與我姊姊大大較力，並且得勝了。」
GEN|30|9|利亞 見自己停了生育，就把她的婢女 悉帕 給 雅各 為妾。
GEN|30|10|利亞 的婢女 悉帕 為 雅各 生了一個兒子。
GEN|30|11|利亞 給他起名叫 迦得 ，說：「真是幸運！」
GEN|30|12|利亞 的婢女 悉帕 又為 雅各 生了第二個兒子。
GEN|30|13|利亞 給他起名叫 亞設 ，說：「我真有福啊，眾女子都要稱我有福。」
GEN|30|14|收割麥子的時候， 呂便 到田裏去，找到曼陀羅草 ，就拿給他的母親 利亞 。 拉結 對 利亞 說：「請你給我一些你兒子的曼陀羅草吧。」
GEN|30|15|利亞 對她說：「你奪走了我的丈夫還是小事嗎？你還要奪取我兒子的曼陀羅草嗎？」 拉結 說：「今夜他可以與你同寢，來交換你兒子的曼陀羅草。」
GEN|30|16|到了晚上， 雅各 從田裏回來， 利亞 出來迎接他，說：「你要與我同寢，因為我真的用我兒子的曼陀羅草把你雇下了。」那一夜， 雅各 就與她同寢。
GEN|30|17|上帝應允了 利亞 ，她就懷孕，為 雅各 生了第五個兒子。
GEN|30|18|利亞 給他起名叫 以薩迦 ，說：「上帝給了我工價，因為我把婢女給了我的丈夫。」
GEN|30|19|利亞 又懷孕，為 雅各 生了第六個兒子。
GEN|30|20|利亞 給他起名叫 西布倫 ，說：「上帝賜給我厚禮了；這次，我丈夫必看重我，因為我為他生了六個兒子。」
GEN|30|21|後來她又生了一個女兒，給她起名叫 底拿 。
GEN|30|22|上帝顧念 拉結 ，應允她，使她能生育。
GEN|30|23|拉結 懷孕生子，說：「上帝除去了我的羞恥。」
GEN|30|24|拉結 就給他起名叫 約瑟 ，說：「願耶和華再增添一個兒子給我。」
GEN|30|25|拉結 生 約瑟 之後， 雅各 對 拉班 說：「請讓我走，回到我的本鄉本土去。
GEN|30|26|請你把我服事你所得的妻子和孩子給我，讓我走吧！我怎樣服事你，你都知道。」
GEN|30|27|拉班 對他說：「願你看得起我，因我占卜得知，耶和華賜福給我是因你的緣故。」
GEN|30|28|又說：「請為我定你的工資，我就給你。」
GEN|30|29|雅各 對他說：「我怎樣服事你，你的牲畜在我這裏變得怎樣，你都知道。
GEN|30|30|我未來以前，你擁有的很少，現在卻已大量增加，因為耶和華隨著我的腳步賜福給你。現在，我到甚麼時候才可以成家立業呢？」
GEN|30|31|拉班 說：「我該給你甚麼呢？」 雅各 說：「你甚麼也不必給我，只要你為我做這件事，我就繼續牧放你的羊群。
GEN|30|32|今天我要走遍你的羊群，把綿羊中凡有點的、有斑的，和小綿羊中凡是黑色的羊；以及山羊中凡有斑的、有點的，都從那裏挑出來，作為我的工資。
GEN|30|33|以後你來當面查看我的工資，任何我這裏的山羊不是有點有斑的，小綿羊不是黑色的，就算是我偷的。這就可以證明我是正直的。」
GEN|30|34|拉班 說：「看哪，就照你所說的做吧。」
GEN|30|35|當日， 拉班 把有紋的、有斑的公山羊，一切有點的、有斑的、有少許白色 的母山羊，以及小綿羊中所有黑色的 ，都挑出來，交在他兒子們的手裏，
GEN|30|36|又使自己和 雅各 相隔三天的路程。 雅各 就牧放 拉班 其餘的羊。
GEN|30|37|雅各 拿楊樹、杏樹、楓樹的嫩枝，把皮剝出白色的條紋，使枝子露出白色來。
GEN|30|38|他把剝了皮的枝子對著羊群，插在羊喝水的水溝和水槽裏。羊來喝水的時候，牠們彼此交配。
GEN|30|39|羊對著枝子交配，就生下有紋的、有點的、有斑的來。
GEN|30|40|雅各 把小綿羊分出來，讓羊對著 拉班 羊群中有紋的和所有黑色的。於是他把自己的羊群分開，不叫牠們和 拉班 的羊混在一起。
GEN|30|41|當肥壯的羊交配的時候， 雅各 就把枝子插在水溝裏，使羊對著枝子交配。
GEN|30|42|可是當瘦弱的羊交配的時候，他就不插枝子。這樣，瘦弱的就歸 拉班 ，肥壯的就歸 雅各 。
GEN|30|43|於是這人極其發達，擁有許多的羊群、奴僕、婢女、駱駝和驢。
GEN|31|1|雅各 聽見 拉班 兒子們的話，說：「 雅各 把我們父親所有的都奪去了！他從我們父親所擁有的獲得這一切的財富。」
GEN|31|2|雅各 見 拉班 的臉色，看哪，待他不如從前了。
GEN|31|3|耶和華對 雅各 說：「你要回你祖先之地，到你本族那裏去，我必與你同在。」
GEN|31|4|雅各 就派人叫 拉結 和 利亞 到田野他的羊群那裏去，
GEN|31|5|對她們說：「我看你們父親待我的臉色不如從前了，但我父親的上帝向來與我同在。
GEN|31|6|你們也知道，我盡了全力服事你們的父親。
GEN|31|7|可是你們的父親欺騙我，十次更改我的工資，但上帝不容許他害我。
GEN|31|8|他若說：『有點的歸給你作工資』，羊群所生的都是有點的；他若說：『有紋的歸給你作工資』，羊群所生的都是有紋的。
GEN|31|9|這樣，上帝把你們父親的牲畜拿來賜給我了。
GEN|31|10|「羊群交配的時候，我在夢中舉目一看，看哪，跳母羊的公羊都是有紋的、有點的、有花斑的。
GEN|31|11|上帝的使者在夢中呼叫我說：『 雅各 。』我說：『我在這裏。』
GEN|31|12|他說：『你舉目觀看，跳母羊的公羊都是有紋的、有點的、有花斑的。 拉班 向你所做的一切，我都看見了。
GEN|31|13|我是 伯特利 的上帝；你曾在那裏用油膏過柱子，向我許過願。現在你起來，離開這地，回你本族之地去吧！』」
GEN|31|14|拉結 和 利亞 回答 雅各 說：「在我們父親家裏還有我們可分得的產業嗎？
GEN|31|15|我們不是被他看作外人嗎？因為他賣了我們，還吞吃了我們的銀錢。
GEN|31|16|上帝從我們父親所拿走的一切財物，都是我們和我們孩子的。現在，凡上帝所吩咐你的，你只管去做吧！」
GEN|31|17|雅各 起來，叫他的孩子和妻子都騎上駱駝，
GEN|31|18|又趕著他一切的牲畜和他所得的一切財物，就是他在 巴旦‧亞蘭 所得的，他擁有的牲畜 ，往 迦南 地他父親 以撒 那裏去了。
GEN|31|19|當時 拉班 去剪羊毛， 拉結 偷了他父親家中的神像。
GEN|31|20|雅各 瞞住 亞蘭 人 拉班 ，不通知他就逃走了。
GEN|31|21|雅各 帶著他所有的逃走了；他起程，渡過 大河 ，面向著 基列山 。
GEN|31|22|到第三天，有人告訴 拉班 ， 雅各 逃跑了。
GEN|31|23|拉班 帶著他的弟兄們去追他，追了七天，就在 基列山 追上了。
GEN|31|24|夜間，上帝來到 亞蘭 人 拉班 那裏，在夢中對他說：「你要小心，不可對 雅各 說好說歹。」
GEN|31|25|拉班 追上 雅各 。 雅各 在山上支搭帳棚； 拉班 和他的弟兄們也在 基列山 上支搭帳棚。
GEN|31|26|拉班 對 雅各 說：「你做的是甚麼事呢？你瞞著我把我的女兒們帶走，好像用刀劍擄去一般。
GEN|31|27|你為甚麼暗暗地逃跑，瞞著我，不通知我一聲，叫我可以歡樂、唱歌、擊鼓、彈琴送你回去呢？
GEN|31|28|為甚麼不容許我與外孫和女兒吻別呢？你現在所做的真是愚蠢！
GEN|31|29|我的手本有能力害你，只是你父親的上帝昨夜對我說：『你要小心，不可對 雅各 說好說歹。』
GEN|31|30|現在你既然這麼想念你的父家，不得不去，為甚麼又偷了我的神明呢？」
GEN|31|31|雅各 回答 拉班 說：「因為我害怕，我想，恐怕你把你的女兒從我這裏奪走。
GEN|31|32|至於你的神明，你若在誰那裏搜出來，就不讓誰活。當著我們弟兄面前，你認一認在我這裏有甚麼東西是你的，你就拿去吧。」原來 雅各 並不知道 拉結 偷了神明。
GEN|31|33|拉班 進了 雅各 、 利亞 ，以及兩個使女的帳棚，卻沒有找到，就從 利亞 的帳棚出來，進入 拉結 的帳棚。
GEN|31|34|拉結 拿了神像，藏在駱駝的鞍子裏，自己坐在上面。 拉班 搜遍了那帳棚，並沒有找到。
GEN|31|35|拉結 對她父親說：「請我主不要生氣，因為我恰有月事，不能在你面前起來。」 拉班 搜尋，卻找不到神像。
GEN|31|36|於是 雅各 發怒，斥責 拉班 。 雅各 對 拉班 說：「我有甚麼過犯，有甚麼罪惡，你竟這樣火速地追我？
GEN|31|37|你搜遍了我一切的物件，你找到甚麼呢？可以放在你我弟兄面前，叫他們在我們兩個之間評評理。
GEN|31|38|我在你那裏這二十年，你的母綿羊、母山羊沒有掉過胎。你羊群中的公綿羊，我沒有吃過；
GEN|31|39|被野獸撕裂的，我沒有帶來給你，是我自己賠償的。無論是白日被偷的，或是黑夜被偷的，你都從我手中索取。
GEN|31|40|我常常白日受盡炎熱，黑夜受盡寒霜，不得合眼入睡。
GEN|31|41|我這二十年在你家裏，為你兩個女兒服事了你十四年，為你的羊群服事了你六年，你卻十次更改我的工資。
GEN|31|42|若不是我父親 以撒 所敬畏的上帝，就是 亞伯拉罕 的上帝與我同在，你如今必定打發我空手而去。上帝看見我的苦情和我手的辛勞，就在昨夜責備了你。」
GEN|31|43|拉班 回答 雅各 說：「這兩個女兒是我的女兒，這些孩子是我的孩子，這些羊群也都是我的羊群；凡你所看見的都是我的。我的女兒和她們所生的孩子，我今日還能對他們做甚麼呢？
GEN|31|44|現在，來吧！讓我和你立約，作你我之間的證據。」
GEN|31|45|雅各 就拿一塊石頭立作柱子，
GEN|31|46|對弟兄們說：「大家來堆積石頭。」他們拿石頭堆成一堆，於是在那裏，在石堆旁邊吃喝。
GEN|31|47|拉班 稱那石堆為 伊迦爾‧撒哈杜他 ， 雅各 卻稱那石堆為 迦累得 。
GEN|31|48|拉班 說：「今日這石堆成為你我之間的證據。」因此這地方名叫 迦累得 ，
GEN|31|49|又叫 米斯巴 ，因為他說：「我們彼此離別以後，願耶和華在你我中間鑒察 。
GEN|31|50|你若苦待我的女兒，或在我的女兒以外另娶妻，雖沒有人在場，你看，有上帝在你我中間作證。」
GEN|31|51|拉班 又對 雅各 說：「看哪，這石堆，看哪，這柱子，是我在你我中間所立的。
GEN|31|52|這石堆是證據，這柱子也是證據。我必不越過這石堆去害你；你也不可越過這石堆和柱子來害我。
GEN|31|53|願 亞伯拉罕 的上帝和 拿鶴 的上帝，就是他們父親的上帝 ，在你我中間判斷。」 雅各 就指著他父親 以撒 所敬畏的上帝起誓，
GEN|31|54|又在山上獻祭，請弟兄們來吃飯。他們吃了飯，就在山上過夜。
GEN|31|55|拉班 清早起來，與他外孫和女兒親吻，為他們祝福，就回到自己的地方去了。
GEN|32|1|雅各 繼續行路，上帝的使者遇見他。
GEN|32|2|雅各 看見他們就說：「這是上帝的軍營。」於是給那地方起名叫 瑪哈念 。
GEN|32|3|雅各 派使者在他前面到 西珥 地，就是 以東 地他哥哥 以掃 那裏。
GEN|32|4|他吩咐他們說：「你們要對我主 以掃 說：『你的僕人 雅各 這樣說：我在 拉班 那裏寄居，延遲到如今。
GEN|32|5|我有牛、驢、羊群、奴僕、婢女，現在派人來報告我主，為了要在你眼前蒙恩。』」
GEN|32|6|使者回到 雅各 那裏，說：「我們到了你哥哥 以掃 那裏。他正迎著你來，並且有四百人和他一起。」
GEN|32|7|雅各 就很懼怕，而且愁煩。他把跟他同行的人和羊群、牛群、駱駝分成兩隊，
GEN|32|8|說：「 以掃 若來擊殺其中一隊，剩下的另一隊還可以逃脫。」
GEN|32|9|雅各 說：「耶和華—我祖父 亞伯拉罕 的上帝，我父親 以撒 的上帝啊，你曾對我說：『回你本地本族去，我要厚待你。』
GEN|32|10|你向僕人所施的一切慈愛和信實，我一點也不配得。我先前只用我的一根杖過這 約旦河 ，如今我卻成了兩隊。
GEN|32|11|求你救我脫離我哥哥的手，脫離 以掃 的手，因為我怕他來殺我，連母親和兒女都不放過。
GEN|32|12|你曾說：『我必定厚待你，使你的後裔如同海邊的沙，多得不可勝數。』」
GEN|32|13|當夜， 雅各 在那裏住宿，就從他手中所擁有的拿禮物要送給他哥哥 以掃 ，
GEN|32|14|就是二百隻母山羊、二十隻公山羊、二百隻母綿羊、二十隻公綿羊、
GEN|32|15|三十匹哺乳的母駱駝和牠們的小駱駝、四十頭母牛、十頭公牛、二十匹母驢和十匹公驢。
GEN|32|16|他把每種牲畜各分一群，交在僕人手中，對僕人說：「你們要在我的前頭過去，使群和群之間保持一段距離」。
GEN|32|17|他又吩咐領頭的人說：「我哥哥 以掃 遇見你的時候，問你說：『你是誰的人？要往哪裏去？你前面這些是誰的？』
GEN|32|18|你就說：『是你僕人 雅各 的，是送給我主 以掃 的禮物。看哪，他自己也在我們後面。』」
GEN|32|19|他又吩咐第二、第三和所有趕畜群的人說：「你們遇見 以掃 的時候要照這樣的話對他說，
GEN|32|20|你們還要說：『看哪，你僕人 雅各 在我們後面。』」因 雅各 說：「我藉著在我前面送去的禮物給他面子，然後再見他的面，或許他會寬容我。」
GEN|32|21|於是禮物在他前面過去了；那夜， 雅各 在營中住宿。
GEN|32|22|他夜間起來，帶著兩個妻子，兩個婢女和十一個孩子，過了 雅博 渡口。
GEN|32|23|他帶著他們，送他們過河，他所有的一切也都過去，
GEN|32|24|只剩下 雅各 一人。有一個人來和他摔跤，直到黎明。
GEN|32|25|那人見自己勝不過他，就摸了他的大腿窩一下。 雅各 的大腿窩就在和那人摔跤的時候扭了。
GEN|32|26|那人說：「天快亮了，讓我走吧！」 雅各 說：「你不給我祝福，我就不讓你走。」
GEN|32|27|那人說：「你叫甚麼名字？」他說：「 雅各 。」
GEN|32|28|那人說：「你的名字不要再叫 雅各 ，要叫 以色列 ，因為你與上帝和人較力，都得勝了。」
GEN|32|29|雅各 問他說：「請告訴我你的名字。」那人說：「何必問我的名字呢？」於是他在那裏為 雅各 祝福。
GEN|32|30|雅各 就給那地方起名叫 毗努伊勒 ，說：「我面對面見了上帝，我的性命仍得保全。」
GEN|32|31|太陽剛出來的時候， 雅各 經過 毗努伊勒 ，他的大腿就瘸了。
GEN|32|32|因此， 以色列 人不吃大腿窩的筋，直到今日，因為那人摸了 雅各 大腿窩的筋。
GEN|33|1|雅各 舉目觀看，看哪， 以掃 來了，有四百人和他一起。 雅各 就把孩子們分開交給 利亞 、 拉結 和兩個婢女。
GEN|33|2|他叫兩個婢女和她們的孩子走在前頭， 利亞 和她的孩子跟在後面，而 拉結 和 約瑟 在最後。
GEN|33|3|他自己卻走到他們前面，一連七次俯伏在地才挨近他哥哥。
GEN|33|4|以掃 跑來迎接他，將他抱住，伏在他的頸項上親他，他們都哭了。
GEN|33|5|以掃 舉目看見婦人和孩子，就說：「這些和你一起的是誰呢？」 雅各 說：「這些孩子是上帝施恩給你僕人的。」
GEN|33|6|於是兩個婢女和她們的孩子前來下拜，
GEN|33|7|利亞 和她的孩子也前來下拜，隨後 約瑟 和 拉結 也前來下拜。
GEN|33|8|以掃 說：「我所遇見的這些畜群是甚麼意思呢？」 雅各 說：「是為了要在我主眼前蒙恩。」
GEN|33|9|以掃 說：「弟弟啊，我的已經夠了，你的你自己留著吧！」
GEN|33|10|雅各 說：「不，我若在你眼前蒙恩，就請你從我手裏收下這禮物；因為我見了你的面，如同見了上帝的面，並且你也寬容了我。
GEN|33|11|請你收下我帶來給你的禮物，因為上帝恩待我，使我一切都充足。」 雅各 再三求他，他才收下。
GEN|33|12|以掃 說：「讓我們起身前行，我和你一起走吧。」
GEN|33|13|雅各 對他說：「我主知道孩子們還年幼嬌嫩，我的牛羊也正在哺乳中，只要催趕一天，群羊都會死了。
GEN|33|14|請我主在僕人前面先走，我要按著在我面前的牲畜和孩子的步伐慢慢前進，直走到 西珥 我主那裏。」
GEN|33|15|以掃 說：「讓我把跟隨我的人留幾個在你這裏。」 雅各 說：「何必這樣呢？只要能在我主眼前蒙恩就夠了。」
GEN|33|16|於是， 以掃 當日起行，回 西珥 去了。
GEN|33|17|雅各 就往 疏割 去，在那裏為自己蓋房屋，又為牲畜搭棚，因此那地方叫 疏割 。
GEN|33|18|雅各 從 巴旦‧亞蘭 平安地回到 迦南 地的 示劍城 ，他在城的前面支搭帳棚。
GEN|33|19|他用一百可錫塔 從 示劍 的父親 哈抹 的眾子手中買了搭帳棚的那塊地。
GEN|33|20|雅各 在那裏築了一座壇，起名叫 伊利‧伊羅伊‧以色列 。
GEN|34|1|利亞 給 雅各 所生的女兒 底拿 出去，要探望那地的女子們。
GEN|34|2|那地的族長 希未 人 哈抹 的兒子 示劍 看見她，就拉住她，與她同寢，玷辱了她。
GEN|34|3|示劍 的心喜歡 雅各 的女兒 底拿 ，愛上這少女，甜言蜜語地安慰她。
GEN|34|4|示劍 對他父親 哈抹 說：「求你為我聘這女孩為妻。」
GEN|34|5|雅各 聽見 示劍 污辱了他的女兒 底拿 。那時他的兒子們正和牲畜在田野， 雅各 就沉默，等他們回來。
GEN|34|6|示劍 的父親 哈抹 出來，到 雅各 那裏，要和他講話。
GEN|34|7|雅各 的兒子們聽見這事，就從田野回來，人人悲憤，十分惱怒，因 示劍 在 以色列 中做了醜事，與 雅各 的女兒同寢，這本是不該做的事。
GEN|34|8|哈抹 和他們談話，說：「我兒子 示劍 的心喜歡你們家的女兒，請你們把她嫁給我的兒子。
GEN|34|9|你們與我們彼此結親；你們可以把你們家的女兒嫁給我們，也可以娶我們家的女兒。
GEN|34|10|你們與我們同住吧！這地都在你們面前，只管在這裏居住，做買賣，置產業。」
GEN|34|11|示劍 對女子的父親和兄弟們說：「願你們看得起我，你們向我要甚麼，我必給你們，
GEN|34|12|無論向我要多貴重的聘金和禮物，我必照你們所說的給你們，只要你們將這少女嫁給我。」
GEN|34|13|雅各 的兒子們因 示劍 污辱了他們的妹妹 底拿 ，就用詭詐的話回答 示劍 和他父親 哈抹 ，
GEN|34|14|對他們說：「我們不能做這樣的事，把我們的妹妹嫁給沒有受割禮的人為妻，因為那是我們的羞恥。
GEN|34|15|惟有一個條件，我們才答應你們，就是你們所有的男丁都要受割禮，和我們一樣，
GEN|34|16|我們就把我們家的女兒嫁給你們，也娶你們家的女兒；我們就與你們同住，大家成為一族人。
GEN|34|17|倘若你們不聽從我們受割禮，我們就帶我們家的女兒走了。」
GEN|34|18|這些話在 哈抹 和他兒子 示劍 的眼中看為美。
GEN|34|19|那年輕人毫不遲延做這事，因為他愛上了 雅各 的女兒；他在他父親家中也是最受人尊重的。
GEN|34|20|哈抹 和他兒子 示劍 到他們的城門口，對城裏的人講說：
GEN|34|21|「這些人對我們友善，不如允許他們在這地居住，做買賣；看哪，這地寬闊，足以容納他們。我們可以娶他們家的女兒，也可以把我們家的女兒嫁給他們。
GEN|34|22|惟有一個條件，這些人才答應和我們同住，成為一族人，就是我們中間所有的男丁都要受割禮，和他們一樣。
GEN|34|23|他們的牲畜、財物和一切的牲口豈不都歸給我們嗎？只要答應他們，他們就與我們同住。」
GEN|34|24|凡從城門出入的人都聽從了 哈抹 和他兒子 示劍 的話。於是，凡從城門出入的男丁都受了割禮。
GEN|34|25|到第三天，他們正疼痛的時候， 雅各 的兩個兒子，就是 底拿 的哥哥 西緬 和 利未 ，各拿刀劍，不動聲色地來到城中，把所有的男丁都殺了，
GEN|34|26|又用刀殺了 哈抹 和他兒子 示劍 ，把 底拿 從 示劍 家裏帶走，就離開了。
GEN|34|27|雅各 的兒子們因為他們的妹妹受污辱，就來到被殺的人那裏，洗劫那城，
GEN|34|28|奪走了他們的羊群、牛群和驢，以及城裏和田間所有的；
GEN|34|29|又俘擄搶劫他們一切的財物、孩童、婦女，以及房屋中所有的。
GEN|34|30|雅各 對 西緬 和 利未 說：「你們連累了我，使我在這地的居民中，就是在 迦南 人和 比利洗 人中壞了名聲。我的人丁稀少，他們必聚集來擊殺我，我和全家的人都要被滅絕。」
GEN|34|31|他們卻說：「他豈可待我們的妹妹如同妓女呢？」
GEN|35|1|上帝對 雅各 說：「起來！上 伯特利 去，住在那裏。在那裏築一座壇給上帝，就是你逃避你哥哥 以掃 的時候向你顯現的上帝。」
GEN|35|2|雅各 就對他家中的人，以及所有和他一起的人說：「除掉你們中間外邦的神明，要自潔，更換衣服。
GEN|35|3|我們要起來，上 伯特利 去，在那裏我要築一座壇給上帝，就是在我遭難的日子應允我，在我行走的路上與我同在的上帝。」
GEN|35|4|他們就把手中所有外邦的神明和自己耳朵上的環子交給 雅各 ； 雅各 把它們埋在 示劍 那裏的橡樹下。
GEN|35|5|他們起行。上帝使周圍城鎮的人都驚恐，就不追趕 雅各 的兒子們了。
GEN|35|6|於是 雅各 和所有與他一起的人到了 迦南 地的 路斯 ，就是 伯特利 。
GEN|35|7|他在那裏築了一座壇，給那地方起名叫 伊勒‧伯特利 ，因為他逃避他哥哥的時候，上帝曾在那裏向他顯現。
GEN|35|8|利百加 的奶媽 底波拉 死了，葬在 伯特利 下邊的橡樹下；那棵樹名叫 亞倫‧巴古 。
GEN|35|9|雅各 從 巴旦‧亞蘭 回來，上帝又向他顯現，賜福給他。
GEN|35|10|上帝對他說：「你的名原是 雅各 ，從今以後不要再叫 雅各 ，你的名要叫 以色列 。」於是，上帝就叫他的名為 以色列 。
GEN|35|11|上帝又對他說：「我是全能的上帝；你要生養眾多，將來有一國和許多的國從你而來，又有許多君王從你生出 。
GEN|35|12|至於我賜給 亞伯拉罕 和 以撒 的地，我必賜給你；我必賜這地給你的後裔。」
GEN|35|13|上帝就從與 雅各 說話的那地方升上去了。
GEN|35|14|雅各 就在上帝與他說話的地方立了一根柱子，就是石柱，在它上面獻澆酒祭，又澆油。
GEN|35|15|雅各 就給上帝與他說話的那地方起名叫 伯特利 。
GEN|35|16|他們從 伯特利 起行，到 以法他 還有一段路程， 拉結 生產，生得十分艱難。
GEN|35|17|她生得十分艱難的時候，接生婆對她說：「不要怕，你又要有一個兒子了。」
GEN|35|18|她快要死，還有一口氣的時候，就給她兒子起名叫 便‧俄尼 ；他父親卻給他起名叫 便雅憫 。
GEN|35|19|拉結 死了，葬在往 以法他 的路旁； 以法他 就是 伯利恆 。
GEN|35|20|雅各 在她的墳上立了一塊碑，就是 拉結 的墓碑，到今日還在。
GEN|35|21|以色列 起行，在 以得臺 的那一邊支搭帳棚。
GEN|35|22|以色列 住在那地的時候， 呂便 去與他父親的妾 辟拉 同寢， 以色列 也聽見了這件事 。 雅各 共有十二個兒子。
GEN|35|23|利亞 的兒子是 雅各 的長子 呂便 ，還有 西緬 、 利未 、 猶大 、 以薩迦 、 西布倫 。
GEN|35|24|拉結 的兒子是 約瑟 、 便雅憫 。
GEN|35|25|拉結 的婢女 辟拉 的兒子是 但 、 拿弗他利 。
GEN|35|26|利亞 的婢女 悉帕 的兒子是 迦得 、 亞設 。這是 雅各 在 巴旦‧亞蘭 所生的兒子。
GEN|35|27|雅各 來到他父親 以撒 那裏，到了 幔利 ， 基列‧亞巴 ，就是 希伯崙 ，是 亞伯拉罕 和 以撒 寄居的地方。
GEN|35|28|以撒 共活了一百八十年。
GEN|35|29|以撒 年紀老邁，安享天年，息勞而終，歸到他祖先 那裏。他兩個兒子 以掃 和 雅各 把他安葬了。
GEN|36|1|這是 以掃 的後代， 以掃 就是 以東 。
GEN|36|2|以掃 娶 迦南 的女子為妻，就是 赫 人 以倫 的女兒 亞大 和 希未 人 祭便 的孫女， 亞拿 的女兒 阿何利巴瑪 ，
GEN|36|3|又娶了 以實瑪利 的女兒， 尼拜約 的妹妹 巴實抹 。
GEN|36|4|亞大 為 以掃 生了 以利法 ； 巴實抹 生了 流珥 ；
GEN|36|5|阿何利巴瑪 生了 耶烏施 、 雅蘭 、 可拉 。這些都是 以掃 的兒子，是在 迦南 地生的。
GEN|36|6|以掃 帶著他的妻子、兒女和家中所有的人，以及他的牛羊、牲畜和一切財物，就是他在 迦南 地所得的，往別處去，離開了他的兄弟 雅各 。
GEN|36|7|因為他們擁有的很多，不能住在一起。因為牲畜的緣故，寄居的地方容不下他們。
GEN|36|8|於是 以掃 住在 西珥山 ； 以掃 就是 以東 。
GEN|36|9|這是 以掃 的後代，他是 西珥山 裏 以東 人的始祖。
GEN|36|10|以掃 子孫的名字如下： 以掃 的妻子 亞大 生 以利法 ； 以掃 的妻子 巴實抹 生 流珥 。
GEN|36|11|以利法 的兒子是 提幔 、 阿抹 、 洗玻 、 迦坦 、 基納斯 。
GEN|36|12|亭納 是 以掃 兒子 以利法 的妾，她為 以利法 生了 亞瑪力 。這是 以掃 的妻子 亞大 的子孫。
GEN|36|13|流珥 的兒子是 拿哈 、 謝拉 、 沙瑪 、 米撒 。這是 以掃 妻子 巴實抹 的子孫。
GEN|36|14|以掃 的妻子 阿何利巴瑪 是 祭便 的孫女， 亞拿 的女兒。她為 以掃 生了 耶烏施 、 雅蘭 、 可拉 。
GEN|36|15|這是 以掃 子孫中作族長的： 以掃 的長子 以利法 的子孫中，有 提幔 族長、 阿抹 族長、 洗玻 族長、 基納斯 族長、
GEN|36|16|可拉 族長、 迦坦 族長、 亞瑪力 族長。這是在 以東 地，從 以利法 所出的族長，是 亞大 的子孫。
GEN|36|17|以掃 的兒子 流珥 的子孫中，有 拿哈 族長、 謝拉 族長、 沙瑪 族長、 米撒 族長。這是在 以東 地，從 流珥 所出的族長，是 以掃 妻子 巴實抹 的子孫。
GEN|36|18|以掃 的妻子 阿何利巴瑪 的子孫中，有 耶烏施 族長、 雅蘭 族長、 可拉 族長。這是從 以掃 的妻子， 亞拿 的女兒 阿何利巴瑪 的子孫中所出的族長。
GEN|36|19|以上的族長都是 以掃 的子孫； 以掃 就是 以東 。
GEN|36|20|這是那地原來的居民， 何利 人 西珥 的子孫： 羅坍 、 朔巴 、 祭便 、 亞拿 、
GEN|36|21|底順 、 以察 、 底珊 。這是在 以東 地，從 何利 人 西珥 子孫中所出的族長。
GEN|36|22|羅坍 的兒子是 何利 、 希幔 ， 羅坍 的妹妹是 亭納 。
GEN|36|23|朔巴 的兒子是 亞勒文 、 瑪拿轄 、 以巴錄 、 示玻 、 阿南 。
GEN|36|24|祭便 的兒子是 愛亞 、 亞拿 ，當時在曠野牧放他父親 祭便 的驢，發現溫泉的就是這 亞拿 。
GEN|36|25|亞拿 的兒子是 底順 ， 亞拿 的女兒是 阿何利巴瑪 。
GEN|36|26|底順 的兒子是 欣但 、 伊是班 、 益蘭 、 基蘭 。
GEN|36|27|以察 的兒子是 辟罕 、 撒番 、 亞干 。
GEN|36|28|底珊 的兒子是 烏斯 、 亞蘭 。
GEN|36|29|這是從 何利 人所出的族長： 羅坍 族長、 朔巴 族長、 祭便 族長、 亞拿 族長、
GEN|36|30|底順 族長、 以察 族長、 底珊 族長。這是從 何利 人所出的族長，都在 西珥 地，按著族長 來分。
GEN|36|31|以色列 未有君王治理之前，這些是在 以東 地作王的。
GEN|36|32|比珥 的兒子 比拉 在 以東 作王，他的城名叫 亭哈巴 。
GEN|36|33|比拉 死了， 波斯拉 人 謝拉 的兒子 約巴 接續他作王。
GEN|36|34|約巴 死了， 提幔 人之地的 戶珊 接續他作王。
GEN|36|35|戶珊 死了， 比達 的兒子 哈達 接續他作王， 哈達 曾在 摩押 地擊敗 米甸 人，他的城名叫 亞未得 。
GEN|36|36|哈達 死了， 瑪士利加 人 桑拉 接續他作王。
GEN|36|37|桑拉 死了， 大河 邊的 利河伯 人 掃羅 接續他作王。
GEN|36|38|掃羅 死了， 亞革波 的兒子 巴勒‧哈南 接續他作王。
GEN|36|39|亞革波 的兒子 巴勒‧哈南 死了， 哈達爾 接續他作王，他的城名叫 巴烏 。他的妻子名叫 米希她別 ，是 米‧薩合 的孫女， 瑪特列 的女兒。
GEN|36|40|這些是 以掃 的族長，按著他們的宗族、住處和名字： 亭納 族長、 亞勒瓦 族長、 耶帖 族長、
GEN|36|41|阿何利巴瑪 族長、 以拉 族長、 比嫩 族長、
GEN|36|42|基納斯 族長、 提幔 族長、 米比薩 族長、
GEN|36|43|瑪基疊 族長、 以蘭 族長。這些是 以東 人在所得為業的地上，按著他們住處的族長。 以掃 是 以東 人的始祖。
GEN|37|1|雅各 住在 迦南 地，就是他父親寄居的地。
GEN|37|2|這是 雅各 的事蹟。 約瑟 十七歲與他哥哥們一同牧羊。他是個少年，與他父親的妾 辟拉 和 悉帕 的兒子們常在一起。 約瑟 把他們的惡行報給父親。
GEN|37|3|以色列 愛 約瑟 過於其他的兒子，因為 約瑟 是他年老生的；他給 約瑟 做了一件長袍 。
GEN|37|4|哥哥們見父親愛 約瑟 過於他們，就恨 約瑟 ，不與他說友善的話。
GEN|37|5|約瑟 做了一個夢，告訴他哥哥們，他們就更加恨他。
GEN|37|6|約瑟 對他們說：「請聽我做的這個夢：
GEN|37|7|看哪，我們在田裏捆禾稼；看哪，我的捆起來站著；看哪，你們的捆圍著我的捆下拜。」
GEN|37|8|他的哥哥們對他說：「難道你真的要作我們的王嗎？難道你真的要統治我們嗎？」他們就因他的夢和他的話更加恨他。
GEN|37|9|後來他又做了另一個夢，告訴他哥哥們說：「看哪，我又做了一個夢；看哪，太陽、月亮和十一顆星都向我下拜。」
GEN|37|10|約瑟 告訴他父親和哥哥們，他父親就責備他說：「你做的這是甚麼夢！難道我和你母親、你的兄弟真的要俯伏在地，來向你下拜嗎？」
GEN|37|11|他的哥哥們都嫉妒他，他父親卻把這事存在心裏。
GEN|37|12|約瑟 的哥哥們到 示劍 去放他們父親的羊。
GEN|37|13|以色列 對 約瑟 說：「你哥哥們不是在 示劍 放羊嗎？來，我派你到他們那裏去。」 約瑟 對他說：「我在這裏。」
GEN|37|14|以色列 對他說：「你去看看你哥哥們是否平安，羊群是否平安，再回來告訴我。」於是他派 約瑟 出 希伯崙谷 ， 約瑟 就往 示劍 去了。
GEN|37|15|有人遇見他，看哪，他在田野走迷了路。那人問他說：「你找甚麼？」
GEN|37|16|他說：「我找我的哥哥們，請告訴我，他們在哪裏放羊。」
GEN|37|17|那人說：「他們已經離開這裏走了，我聽見他們說：『我們往 多坍 去。』」 約瑟 就去追哥哥們，在 多坍 找到了他們。
GEN|37|18|他們遠遠看見他，趁他還沒有走近他們，就圖謀要殺死他。
GEN|37|19|他們彼此說：「看哪！那做夢的來了。
GEN|37|20|現在，來吧！我們把他殺了，丟在一個坑裏，就說有惡獸把他吃了。我們且看他的夢將來怎麼樣。」
GEN|37|21|呂便 聽見了，要救 約瑟 脫離他們的手，說：「我們不可害他的性命」；
GEN|37|22|呂便 又對他們說：「不可流他的血，可以把他丟在這曠野的坑裏，不可下手害他。」 呂便 要救他脫離他們的手，把他還給他父親。
GEN|37|23|約瑟 到了他哥哥們那裏，他們就剝去他的外衣，就是他身上那件長袍。
GEN|37|24|他們抓住他，把他丟在坑裏。那坑是空的，裏頭沒有水。
GEN|37|25|他們坐下吃飯，舉目觀看，看哪，有一群 以實瑪利 人從 基列 來，用駱駝馱著香料、乳香、沒藥，要帶下 埃及 去。
GEN|37|26|猶大 對他的兄弟們說：「我們殺我們的弟弟，遮掩他的血有甚麼好處呢？
GEN|37|27|來，我們把他賣給 以實瑪利 人，不要下手害他，因為他是我們的弟弟，我們的骨肉。」他的兄弟們就聽從了他。
GEN|37|28|那時，有些 米甸 的商人從那裏經過，就把 約瑟 從坑裏拉上來。他們以二十塊銀子把 約瑟 賣給 以實瑪利 人，他們就把 約瑟 帶到 埃及 去了。
GEN|37|29|呂便 回到坑旁，看哪， 約瑟 不在坑裏，就撕裂自己的衣服，
GEN|37|30|回到他兄弟們那裏，說：「孩子不在了。我往哪裏去才好呢？」
GEN|37|31|於是，他們宰了一隻公山羊，拿了 約瑟 的那件外衣染上了血，
GEN|37|32|派人把長袍送到他們的父親那裏，說：「我們發現這個， 請認一認，是不是你兒子的外衣？」
GEN|37|33|他認出來，就說：「這是我兒子的外衣，惡獸把他吃了， 約瑟 一定被撕碎了！」
GEN|37|34|雅各 就撕裂衣服，腰間圍上麻布，為他兒子哀傷了多日。
GEN|37|35|他的兒女都起來安慰他，他卻不肯受安慰，說：「我必哀傷著下陰間，到我兒子那裏。」 約瑟 的父親就為他哀哭。
GEN|37|36|米甸 人把 約瑟 賣到 埃及 ，給法老的官員，就是護衛長 波提乏 。
GEN|38|1|那時， 猶大 離開他兄弟們下去，到一個名叫 希拉 的 亞杜蘭 人的家附近支搭帳棚。
GEN|38|2|猶大 在那裏看見一個名叫 拔．書亞 的 迦南 女子，就娶她為妻，與她同房，
GEN|38|3|她就懷孕生了兒子， 猶大 給他起名叫 珥 。
GEN|38|4|她又懷孕生了兒子，給他起名叫 俄南 。
GEN|38|5|她又再生了兒子，給他起名叫 示拉 。她生 示拉 的時候， 猶大 正在 基悉 。
GEN|38|6|猶大 為長子 珥 娶妻，名叫 她瑪 。
GEN|38|7|猶大 的長子 珥 在耶和華眼中看為惡，耶和華就殺死了他。
GEN|38|8|猶大 對 俄南 說：「你當與你哥哥的妻子同房，向她盡你的本分，為你哥哥生子立後。」
GEN|38|9|俄南 知道如果與嫂嫂同房，所生的孩子不屬於自己，就洩在地上，不為哥哥生子立後。
GEN|38|10|俄南 所做的在耶和華眼中看為惡，耶和華也殺死了他。
GEN|38|11|猶大 對他媳婦 她瑪 說：「你去住在你父親家裏守寡，等我兒子 示拉 長大。」因為他說：「恐怕 示拉 也像兩個哥哥一樣死去。」 她瑪 就去，住在她父親家裏。
GEN|38|12|過了一段很長的日子， 猶大 的妻子， 書亞 的女兒死了。 猶大 受到了安慰，就和他朋友 亞杜蘭 人 希拉 上 亭拿 去，到他的剪羊毛的人那裏。
GEN|38|13|有人告訴 她瑪 說：「看哪，你的公公上 亭拿 剪羊毛去了。」
GEN|38|14|她瑪 見 示拉 已經長大，卻還沒有娶她為妻，就脫去她寡婦的衣裳，用面紗蒙著，蓋住自己，坐在往 亭拿 的路上， 伊拿印 城門口。
GEN|38|15|猶大 看見她，以為是妓女，因為她蒙著臉。
GEN|38|16|猶大 就轉到路邊她那裏，說：「來吧！讓我與你同寢。」他並不知道她就是他的媳婦。 她瑪 說：「你要與我同寢，把甚麼給我呢？」
GEN|38|17|猶大 說：「我從羊群裏取一隻小山羊，派人送來給你。」 她瑪 說：「在未送之前，你能給我一個信物嗎？」
GEN|38|18|他說：「我給你甚麼信物呢？」 她瑪 說：「你的印、你的帶子 和你手裏的杖。」於是 猶大 給了她，與她同寢，她就從 猶大 懷了孕。
GEN|38|19|她瑪 起來走了，除去面紗，照常穿上寡婦的衣裳。
GEN|38|20|猶大 託他朋友 亞杜蘭 人送一隻小山羊去，要從那女人手裏取回信物，卻找不到她。
GEN|38|21|他問那地方的人說：「 伊拿印 路旁的神廟娼妓在哪裏？」他們說：「這裏沒有神廟娼妓。」
GEN|38|22|他回到 猶大 那裏說：「我找不到她，並且那地方的人說：『這裏沒有神廟娼妓。』」
GEN|38|23|猶大 說：「讓她拿去吧，免得我們被人譏笑。看哪，我把這小山羊送去了，可是你找不到她。」
GEN|38|24|大約過了三個月，有人告訴 猶大 說：「你的媳婦 她瑪 行淫，並且，看哪，她因行淫而懷了孕。」 猶大 說：「拉她出來，把她燒了！」
GEN|38|25|她瑪 被拉出來的時候，就派人到她公公那裏，對他說：「這些東西是誰的，我就是從誰懷了孕。」她又說：「請你認一認，這印、這帶子和這杖是誰的？」
GEN|38|26|猶大 承認說：「她比我更有理，因為我沒有把她給我的兒子 示拉 。」 猶大 再也不跟她同寢。
GEN|38|27|她瑪 生產的時候到了，看哪，腹裏懷的是雙胞胎。
GEN|38|28|生產的時候，一個孩子伸出手來；接生婆拿紅線綁在他手上，說：「這是頭生的。」
GEN|38|29|這孩子把手收回去，看哪，他哥哥生出來了；接生婆說：「你竟然為自己衝出一個裂縫！」於是，他的名字叫 法勒斯 。
GEN|38|30|後來，那手上有紅線的兄弟也生出來，他的名字叫 謝拉 。
GEN|39|1|約瑟 被帶下 埃及 去。有一個 埃及 人 波提乏 ，是法老的官員，是護衛長，他從那些帶 約瑟 下來的 以實瑪利 人手中把 約瑟 買了去。
GEN|39|2|約瑟 在他 埃及 主人的家中，耶和華與他同在，他是一個通達的人。
GEN|39|3|他主人見耶和華與他同在，又見耶和華使他手裏所辦的事都順利，
GEN|39|4|約瑟 就在主人眼前蒙恩，伺候他主人，主人派他管理家務，把一切所有的都交在他手裏。
GEN|39|5|自從主人派 約瑟 管理家務和他一切所有的，耶和華就因 約瑟 的緣故賜福給那 埃及 人的家；凡家裏和田間一切所有的，都蒙耶和華賜福。
GEN|39|6|波提乏 把他一切所有的都交在 約瑟 手中，除了自己所吃的食物，其他的事一概不知。 約瑟 英俊健美。
GEN|39|7|這些事以後， 約瑟 主人的妻子以目送情給 約瑟 ，說：「你與我同寢吧！」
GEN|39|8|約瑟 拒絕，對他主人的妻子說：「看哪，一切家務我主人一概不知，他把所有的都交在我手裏。
GEN|39|9|在這家裏沒有人比我更大，除你以外，他也沒有留下一樣不交給我，因為你是他的妻子。我怎能行這麼大的惡，得罪上帝呢？」
GEN|39|10|她天天這樣對 約瑟 說， 約瑟 卻不聽從她，不與她同寢，也不和她在一起。
GEN|39|11|有一天， 約瑟 進屋裏去辦事，家裏沒有一個人在那屋子裏，
GEN|39|12|婦人就拉住他的衣服，說：「你與我同寢吧！」 約瑟 把衣服留在她手裏，逃出外面去了。
GEN|39|13|婦人看見 約瑟 把衣服留在她手裏逃到外面，
GEN|39|14|就叫了家裏的人來，對他們說：「看，他帶了一個 希伯來 人到我們這裏戲弄我們。他到我這裏來，要與我同寢，我就大聲喊叫。
GEN|39|15|他聽見我放聲大喊，就把他的衣服留在我這裏，逃出外面去了。」
GEN|39|16|婦人把 約瑟 的衣服放在身邊，直到他主人回家，
GEN|39|17|就用這樣的話對他說：「你帶到我們這裏來的那 希伯來 僕人進來要調戲我，
GEN|39|18|我放聲大喊，他就把衣服留在我身邊，逃到外面。」
GEN|39|19|主人聽見他妻子對他說的話，說：「你的僕人就是這樣對待我」，就非常生氣。
GEN|39|20|約瑟 的主人把他抓起來，關在監獄裏，就是王的囚犯被關的地方。於是 約瑟 在那裏坐牢。
GEN|39|21|但耶和華與 約瑟 同在，向他施恩，使他在監獄長的眼前蒙恩。
GEN|39|22|監獄長就把監獄裏所有的囚犯都交在 約瑟 手下；在那裏的一切事都由他處理。
GEN|39|23|任何交在 約瑟 手中的事，監獄長一概不察，因為耶和華與 約瑟 同在，耶和華使他所做的都順利。
GEN|40|1|這些事以後， 埃及 王的司酒長和司膳長得罪了他們的主 埃及 王。
GEN|40|2|法老就對司酒長和司膳長兩個官員發怒，
GEN|40|3|把他們關在護衛長府內的監獄裏，就是 約瑟 被囚的地方。
GEN|40|4|護衛長把他們交給 約瑟 ， 約瑟 就伺候他們。他們被關了一段日子。
GEN|40|5|關在監獄裏的這兩個人，就是 埃及 王的司酒長和司膳長，在同一個晚上各自做了一個夢，每個夢都有自己的解釋。
GEN|40|6|到了早晨， 約瑟 來到他們那裏看他們，看哪，他們很憂愁。
GEN|40|7|他就問一同關在他主人府內法老的官員，說：「你們今日為甚麼面帶愁容呢？」
GEN|40|8|他們對他說：「我們各自做了一個夢，卻沒有人能講解。」 約瑟 對他們說：「解夢不是出於上帝嗎？請你們把夢告訴我。」
GEN|40|9|司酒長就把夢告訴 約瑟 ，對他說：「在我的夢中，看哪，有一棵葡萄樹在我面前，
GEN|40|10|樹上有三根枝子。枝子發了芽，開了花，結出串串成熟的葡萄。
GEN|40|11|法老的杯在我手中，我就拿葡萄擠在法老的杯裏，把杯遞到他手中。」
GEN|40|12|約瑟 對他說：「夢的解釋是這樣：三根枝子就是三天；
GEN|40|13|三天之內，法老要讓你抬起頭來，叫你官復原職。你仍要遞杯在法老的手中，像先前作他的司酒長一樣。
GEN|40|14|但你得福的時候，請你記得我，向我施慈愛，在法老面前提起我，救我出這監牢。
GEN|40|15|我實在是從 希伯來 人之地被拐來的，我在這裏也沒有做過甚麼，好叫他們把我關在牢裏。」
GEN|40|16|司膳長見夢解得好，就對 約瑟 說：「在我夢中，看哪，我頭上頂著三個裝餅的籃子；
GEN|40|17|最上面的籃子裏有為法老烤的各樣食物，有飛鳥來吃我頭上籃子裏的食物。」
GEN|40|18|約瑟 說：「夢的解釋是這樣：三個籃子就是三天；
GEN|40|19|三天之內，法老要讓你抬起頭來，身首異處，把你掛在木架上，必有飛鳥來吃你身上的肉。」
GEN|40|20|到了第三天，正是法老的生日，他為眾臣僕擺設宴席，使司酒長和司膳長從眾臣僕中抬起頭來，
GEN|40|21|讓司酒長官復原職，仍舊遞杯在法老手中，
GEN|40|22|卻把司膳長掛起來，正如 約瑟 向他們所講解的。
GEN|40|23|然而，司酒長不記得 約瑟 ，竟忘了他。
GEN|41|1|過了兩年，法老做夢，看哪，自己站在 尼羅河 邊，
GEN|41|2|看哪，有七頭母牛從 尼羅河 裏上來，長相俊美，肌肉肥壯，在蘆葦中吃草。
GEN|41|3|看哪，隨後又有七頭母牛從 尼羅河 裏上來，長相醜陋，肌肉乾瘦，與那七頭母牛一同站在河邊。
GEN|41|4|這長相醜陋，肌肉乾瘦的七頭母牛吃了那長相俊美又肥壯的七頭母牛。法老就醒了。
GEN|41|5|他又睡著，第二次做夢，看哪，一株麥桿長了七個穗子，又肥大又佳美，
GEN|41|6|看哪，隨後又長出七個穗子，又細弱又被東風吹焦了。
GEN|41|7|這細弱的穗子吞了那七個又肥大又飽滿的穗子。法老醒了，看哪，是個夢。
GEN|41|8|到了早晨，法老心裏不安，就派人把 埃及 所有的術士和智慧人都召來。法老把所做的夢告訴他們，但是沒有人能為法老解夢。
GEN|41|9|那時司酒長對法老說：「我今日想起我的罪來。
GEN|41|10|從前法老對臣僕發怒，把我和司膳長關在護衛長府內的監牢裏。
GEN|41|11|我們兩人在同一晚上各做一夢，每個夢都有各自的解釋。
GEN|41|12|同我們在一起有一個 希伯來 的年輕人，是護衛長的僕人。我們告訴他，他就為我們解夢，照著各人的夢講解。
GEN|41|13|後來事情正如他給我們講解的實現了，我官復原職，司膳長被掛起來了。」
GEN|41|14|於是法老派人去召 約瑟 ，他們就急忙把他從牢裏提出來。他就剃頭刮臉，換衣服，進到法老面前。
GEN|41|15|法老對 約瑟 說：「我做了一個夢，沒有人能講解。我聽人說，你聽了夢就能講解。」
GEN|41|16|約瑟 回答法老說：「這不在乎我。上帝必應允法老平安。」
GEN|41|17|法老對 約瑟 說：「在我的夢中，看哪，我站在 尼羅河 邊，
GEN|41|18|看哪，有七頭母牛從 尼羅河 裏上來，肌肉肥壯，外形俊美，在蘆葦中吃草。
GEN|41|19|看哪，隨後又有七頭母牛上來，虛弱，外形很醜陋，肌肉又乾瘦，在 埃及 全地，我沒有見過這樣醜陋的牛。
GEN|41|20|這乾瘦又醜陋的母牛吃了那先前的七頭肥母牛，
GEN|41|21|進了肚子以後卻看不出已經進了肚子，那醜陋的長相仍舊和先前一樣。我就醒了。
GEN|41|22|我又在夢中觀看，看哪，一株麥桿長了七個穗子，又飽滿又佳美，
GEN|41|23|看哪，隨後又長出七個穗子，枯槁，細弱，又被東風吹焦了。
GEN|41|24|這些細弱的穗子吞了那七個佳美的穗子。我告訴術士，卻沒有人能為我講解。」
GEN|41|25|約瑟 對法老說：「法老的夢是同一個。上帝已把要做的事指示法老了。
GEN|41|26|七頭好母牛是七年，七個佳美的穗子也是七年，這是同一個夢。
GEN|41|27|那隨後上來的七頭乾瘦又醜陋的母牛是七年；那七個空心，被東風吹焦的穗子也一樣，都是七個荒年。
GEN|41|28|這就是我對法老所說，上帝已把要做的事顯明給法老了。
GEN|41|29|看哪，必有七個大豐年來到 埃及 全地，
GEN|41|30|隨後又有七個荒年，甚至 埃及 地的人都忘了先前的豐收，這地必被饑荒所滅。
GEN|41|31|因為那後來的饑荒非常嚴重，就不覺得這地先前有豐收。
GEN|41|32|至於法老兩次做夢，是因為上帝已經確定這事，上帝必速速成就。
GEN|41|33|現在，請法老選一個聰明又有智慧的人，委派他治理 埃及 地。
GEN|41|34|請法老這樣做，委派官員治理這地，在七個豐年的期間，徵收 埃及 地出產的五分之一，
GEN|41|35|叫他們聚集未來豐年一切的糧食，積存五穀歸在法老的手下作糧食，儲藏在各城裏。
GEN|41|36|這糧食可以為這地作儲備，為了 埃及 地要來的七個荒年，免得這地被饑荒所滅。」
GEN|41|37|這事在法老和他眾臣僕眼中都覺得好。
GEN|41|38|法老對臣僕說：「像這樣的人，有上帝的靈在他裏面，我們豈能找得著呢？」
GEN|41|39|法老對 約瑟 說：「上帝既指示你這一切事，就沒有人像你這樣聰明又有智慧。
GEN|41|40|你可以治理我的家；我的百姓都必服從你口中的命令。惟獨在寶座上，我比你大。」
GEN|41|41|法老又對 約瑟 說：「看，我委派你治理 埃及 全地。」
GEN|41|42|法老就脫下手上帶印的戒指，戴在 約瑟 的手上，給他穿上細麻衣，把金鏈戴在他的頸項上，
GEN|41|43|又給 約瑟 坐他的副座車，在他前面有人呼叫說：「跪下 。」於是，法老委派他治理 埃及 全地。
GEN|41|44|法老對 約瑟 說：「我是法老，若沒有你的命令， 埃及 全地的人都不可擅自辦事 。」
GEN|41|45|法老給 約瑟 起名叫 撒發那特‧巴內亞 ，又將 安城 的祭司 波提‧非拉 的女兒 亞西納 給他為妻。 約瑟 就出去治理 埃及 地。
GEN|41|46|約瑟 在 埃及 王法老面前侍立的時候年三十歲。 約瑟 從法老面前出去，巡行 埃及 全地。
GEN|41|47|七個豐年之內，地的出產極其豐盛 ，
GEN|41|48|約瑟 聚集 埃及 地七年一切的糧食，把糧食積存在各城裏，就是把各城周圍田地的糧食都積存在該城裏。
GEN|41|49|約瑟 積存的五穀很多，如同海邊的沙，無法計算，數也數不清。
GEN|41|50|荒年未到以前， 安城 的祭司 波提‧非拉 的女兒 亞西納 為 約瑟 生了兩個兒子。
GEN|41|51|約瑟 給長子起名叫 瑪拿西 ，因為他說：「上帝使我忘了一切的困苦和我父的全家。」
GEN|41|52|他給次子起名叫 以法蓮 ，因為他說：「上帝使我在受苦的地方興盛。」
GEN|41|53|埃及 地的七個豐年一過，
GEN|41|54|七個荒年就來了，正如 約瑟 所說的。各地都有饑荒，惟獨 埃及 全地有糧食。
GEN|41|55|等到 埃及 全地也有了饑荒，眾百姓就向法老哀求糧食。法老對所有的 埃及 人說：「你們到 約瑟 那裏去，凡他所說的，你們都要做。」
GEN|41|56|當時饑荒遍滿了全地， 約瑟 就開了各處的糧倉 ，賣糧食給 埃及 人。 埃及 地的饑荒非常嚴重。
GEN|41|57|各地的人都去 埃及 ，到 約瑟 那裏買糧食，因為全地的饑荒非常嚴重。
GEN|42|1|雅各 見 埃及 有糧，就對兒子們說：「你們為甚麼彼此對看呢？」
GEN|42|2|他又說：「看哪，我聽見 埃及 有糧，你們可以下到那裏，從那裏為我們買些糧來，我們就可以存活，不至於死。」
GEN|42|3|於是， 約瑟 的十個哥哥都下去，到 埃及 買糧食。
GEN|42|4|至於 約瑟 的弟弟 便雅憫 ， 雅各 沒有派他和哥哥們同去，因為 雅各 說：「恐怕他遭難。」
GEN|42|5|以色列 的兒子們來了，在前來的人當中，為要買糧食，因為 迦南 地也有饑荒。
GEN|42|6|當時在 埃及 地掌權的人是 約瑟 ，賣糧給各地眾百姓的就是他。 約瑟 的哥哥們來了，臉伏於地，向他下拜。
GEN|42|7|約瑟 看見他哥哥們，就認出他們，卻對他們裝作陌生人，向他們說嚴厲的話，對他們說：「你們從哪裏來？」他們說：「我們從 迦南 地來買糧。」
GEN|42|8|約瑟 認得他哥哥們，他們卻不認得他。
GEN|42|9|約瑟 想起從前所做的那兩個夢，就對他們說：「你們是奸細，你們來是要窺探這地的虛實。」
GEN|42|10|他們對他說：「我主啊，不是的，僕人們是來買糧的。
GEN|42|11|我們都是同一個人的兒子，我們是誠實的人。僕人們並不是奸細。」
GEN|42|12|約瑟 對他們說：「不，你們一定是窺探這地的虛實來的。」
GEN|42|13|他們說：「僕人們本是兄弟十二人，我們都是 迦南 地同一個人的兒子。看哪，最小的今日在我們父親那裏，有一個不在了。」
GEN|42|14|約瑟 對他們說：「我剛才對你們說過了，你們是奸細！
GEN|42|15|我指著法老的性命起誓，若是你們最小的弟弟不到這裏來，你們就不可以離開這裏；這樣你們就可以證實自己了。
GEN|42|16|要派你們當中的一個人去，把你們的弟弟帶來。至於你們，都要關在這裏，好證實你們的話是不是真的。若不是，我指著法老的性命起誓，你們一定是奸細。」
GEN|42|17|於是 約瑟 把他們一起都關在監裏三天。
GEN|42|18|第三天， 約瑟 對他們說：「我是敬畏上帝的，你們這麼做就可以活。
GEN|42|19|如果你們是誠實的人，留你們兄弟中的一個關在監牢裏，你們帶糧食回去，救你們家的饑荒，
GEN|42|20|再把你們最小的弟弟帶到我這裏來。如此，你們的話就是真的了，你們也不至於死。」他們就照樣做了。
GEN|42|21|他們彼此說：「我們在弟弟身上實在犯了罪。他哀求我們的時候，我們看見他的痛苦，卻不肯聽，所以這場苦難臨到我們。」
GEN|42|22|呂便 回答他們說：「我不是對你們說過，不可傷害那孩子嗎？只是你們不肯聽，看哪，他的血在追討了。」
GEN|42|23|他們不知道 約瑟 在聽，因為在他們之間有傳譯官。
GEN|42|24|約瑟 轉身離開他們，哭了一場，又回來對他們說話，就從他們中間抓了 西緬 ，在他們眼前捆綁他。
GEN|42|25|約瑟 吩咐人把他們的器皿裝滿糧食，把各人的銀子退還在各人的袋裏，又給他們路上需用的食物。人就為他們這樣做了。
GEN|42|26|他們把糧食馱在驢上，離開那裏去了。
GEN|42|27|到了住宿的地方，有一個人打開袋子，要拿飼料餵驢，就看見自己的銀子，看哪，仍在袋口上。
GEN|42|28|他對兄弟們說：「我的銀子退回來了，看哪，還在我袋子裏！」他們戰戰兢兢，心都快跳出來了，彼此說：「上帝向我們做的是甚麼呢？」
GEN|42|29|他們來到 迦南 地他們的父親 雅各 那裏，把所遭遇的事都告訴他，說：
GEN|42|30|「那地的主對我們說嚴厲的話，把我們當作窺探那地的奸細。
GEN|42|31|我們對他說：『我們是誠實的人，並不是奸細。
GEN|42|32|我們本是兄弟十二人，都是同一個父親的兒子，有一個不在了，最小的今日和我們父親在 迦南 地。』
GEN|42|33|那地的主對我們說：『只有這樣我才知道你們是誠實的人：留你們兄弟中的一個在我這裏，你們帶糧食回去，救你們家的饑荒，
GEN|42|34|再把你們最小的弟弟帶到我這裏來，我就知道你們不是奸細，是誠實的人。然後，我就把你們的兄弟交還你們，你們也可以在此地做買賣。』」
GEN|42|35|後來他們倒空袋子，看哪，各人的銀囊都在袋子裏。他們和父親看見銀囊就都害怕。
GEN|42|36|他們的父親 雅各 對他們說：「你們害我喪失了我的兒子： 約瑟 不在了， 西緬 也不在了，你們還要帶走 便雅憫 ！這些事都臨到我身上了。」
GEN|42|37|呂便 對他父親說：「我若不帶他回來給你，你可以殺我的兩個兒子。只管把他交在我手裏，我必帶他回來給你。」
GEN|42|38|雅各 說：「我的兒子不可與你們一同下去。他哥哥死了，只剩下他。他若在你們行走的路上遭難，你們就害我白髮蒼蒼、悲悲慘慘下陰間去了。」
GEN|43|1|那地的饑荒非常嚴重。
GEN|43|2|他們從 埃及 帶來的糧食吃完了，父親對他們說：「你們再去給我們買些糧來。」
GEN|43|3|猶大 對他說：「那人嚴厲地警告我們說：『你們的弟弟若不和你們同來，你們就不要來見我的面。』
GEN|43|4|你若派我們的弟弟跟我們同去，我們就下去給你買糧；
GEN|43|5|你若不派他去，我們就不下去，因為那人對我們說：『你們的弟弟若不和你們同來，你們就不要來見我的面。』」
GEN|43|6|以色列 說：「你們為甚麼這樣害我，告訴那人你們還有弟弟呢？」
GEN|43|7|他們說：「那人詳細問到我們和我們的家人，說：『你們的父親還在嗎？你們還有兄弟嗎？』我們就按著他的這些話告訴他，我們怎麼知道他會說：『把你們的弟弟帶下來』呢？」
GEN|43|8|猶大 又對他父親 以色列 說：「請派這年輕人和我同去，我們就動身前去，好叫我們和你，以及我們的孩子都得存活，不至於死。
GEN|43|9|我為他擔保，你可以從我手中要人，我若不帶他回來交在你面前，我就對你永遠擔當這罪。
GEN|43|10|我們若沒有耽擱，現在第二趟都回來了。」
GEN|43|11|父親 以色列 對他們說：「如果必須如此，你們要這樣做：把本地土產中最好的乳香、蜂蜜、香料、沒藥、堅果、杏仁各取一點，放在器皿裏，帶下去送給那人作禮物。
GEN|43|12|手裏要帶雙倍的銀子，把退還在你們袋口的銀子親手帶回去；或許那是個失誤。
GEN|43|13|帶著你們的弟弟，動身再去見那人。
GEN|43|14|願全能的上帝使你們在那人面前蒙憐憫，放你們另一個兄弟和 便雅憫 回來。我若要失喪兒子，就喪了吧！」
GEN|43|15|於是，他們拿著那些禮物，手裏也帶雙倍的銀子，並且帶著 便雅憫 ，動身下到 埃及 ，站在 約瑟 面前。
GEN|43|16|約瑟 見 便雅憫 和他們同來，就對管家說：「把這些人領到屋裏。要宰殺牲畜，預備宴席，因為中午這些人要跟我吃飯。」
GEN|43|17|那人就照 約瑟 所說的去做，領他們進 約瑟 的屋裏。
GEN|43|18|這些人因為被領到 約瑟 的屋裏，就害怕，說：「領我們到這裏來，必是因為當初退還在我們袋裏的銀子，要設計害我們，抓我們去當奴隸，搶奪我們的驢。」
GEN|43|19|他們就挨近 約瑟 的管家，在屋子門口和他說話，
GEN|43|20|說：「我主啊，求求你，我們當初下來，真的是要買糧食。
GEN|43|21|後來到了住宿的地方，我們打開袋子，看哪，各人的銀子還在自己的袋口上，銀子的分量一點不少。現在我們親手把它帶回來，
GEN|43|22|我們手裏又帶了另外的銀子來買糧食。我們不知道是誰把銀子放在我們袋裏的。」
GEN|43|23|他說：「你們平安！不要害怕，是你們的上帝和你們父親的上帝把財寶放在你們的袋裏。你們的銀子，我已經收了。」他就把 西緬 帶出來，交給他們。
GEN|43|24|那人領這些人進 約瑟 的屋裏，給他們水洗腳，又給他們飼料餵驢。
GEN|43|25|他們預備好禮物，等候 約瑟 中午來，因為他們聽說他們要在那裏吃飯。
GEN|43|26|約瑟 來到家裏，他們就把手中的禮物拿進屋裏給他，俯伏在地，向他下拜。
GEN|43|27|約瑟 問他們安，又說：「你們的父親，就是你們所說的那位老人家平安嗎？他還在嗎？」
GEN|43|28|他們說：「你僕人，我們的父親平安，他還在。」於是他們低頭下拜。
GEN|43|29|約瑟 舉目看見他同母的弟弟 便雅憫 ，就說：「你們向我所說那最小的弟弟就是這位嗎？」又說：「我兒啊，願上帝賜恩給你！」
GEN|43|30|約瑟 愛弟之情激動，就急忙找個地方去哭。他進入自己的房間，哭了一場。
GEN|43|31|他洗了臉出來，勉強忍住，就說：「開飯吧！」
GEN|43|32|他們為 約瑟 單獨擺了一席，為那些人又擺了一席，也為和 約瑟 同吃飯的 埃及 人另擺了一席，因為 埃及 人不和 希伯來 人一同吃飯；那是 埃及 人所厭惡的。
GEN|43|33|兄弟們被安排在 約瑟 面前坐席，都按著長幼的次序，這些人彼此感到詫異。
GEN|43|34|約瑟 把他面前的食物分給他們，但 便雅憫 所得的比別人多五倍。他們就喝酒，和 約瑟 一同暢飲。
GEN|44|1|約瑟 吩咐管家說：「按照他們的驢子所能馱的，把這些人的袋子裝滿糧食，再把各人的銀子放在各人的袋口上，
GEN|44|2|我的杯，就是那個銀杯，要和買糧的銀子一同放在最年輕的那個人的袋口上。」管家就照 約瑟 所說的話去做了。
GEN|44|3|天一亮，這些人和他們的驢子就被送走了。
GEN|44|4|他們出城走了不遠， 約瑟 對管家說：「起來，去追那些人，追上了就對他們說：『你們為甚麼以惡報善呢？
GEN|44|5|這不是我主人用來飲酒，確實用它來占卜的嗎？你們這麼做是不對的！』」
GEN|44|6|管家追上他們，把這些話對他們說了。
GEN|44|7|他們對他說：「我主為甚麼說這樣的話呢？你僕人們絕不會做這樣的事。
GEN|44|8|看哪，我們從前在袋口上發現的銀子，尚且從 迦南 地帶來還你，我們又怎麼會從你主人家裏偷竊金銀呢？
GEN|44|9|你僕人中無論在誰那裏找到杯子，就叫他死，我們也要作我主的奴隸。」
GEN|44|10|管家說：「現在就照你們的話做吧！在誰那裏找到杯子，誰就作我的奴隸，其餘的人都沒有罪。」
GEN|44|11|於是他們各人急忙把袋子卸在地上，各人打開自己的袋子。
GEN|44|12|管家就搜查，從年長的開始到年幼的為止，那杯竟在 便雅憫 的袋子裏找到了。
GEN|44|13|他們就撕裂衣服，各人把馱子抬在驢上，回城去了。
GEN|44|14|猶大 和他兄弟們來到 約瑟 的屋裏， 約瑟 還在那裏，他們就在他面前俯伏於地。
GEN|44|15|約瑟 對他們說：「你們做的是甚麼事呢？你們豈不知像我這樣的人必懂得占卜嗎？」
GEN|44|16|猶大 說：「我們對我主能說甚麼呢？還有甚麼話可說呢？我們還能為自己表白嗎？上帝已經查出你僕人的罪孽了。看哪，我們與那在他手中找到杯子的人都是我主的奴隸。」
GEN|44|17|約瑟 說：「我絕不能做這樣的事！誰的手中找到杯子，誰就作我的奴隸。至於你們，可以平平安安上到你們父親那裏去。」
GEN|44|18|猶大 挨近他，說：「我主啊，求求你，讓僕人說一句話給我主聽，不要向僕人發烈怒，因為你如同法老一樣。
GEN|44|19|我主曾問僕人們說：『你們有父親、兄弟沒有？』
GEN|44|20|我們對我主說：『我們有父親，他已經年老，還有他老年所生的一個小兒子。他哥哥死了，他的母親只剩下他一個孩子，父親也疼愛他。』
GEN|44|21|你對僕人說：『把他帶下到我這裏來，讓我親眼看看他。』
GEN|44|22|我們對我主說：『這年輕人不能離開他父親，若是離開，父親就會死。』
GEN|44|23|你對僕人說：『你們最小的弟弟若不和你們一同下來，你們就不要來見我的面。』
GEN|44|24|我們上到你僕人，我們父親那裏，就把我主的話告訴了他。
GEN|44|25|後來，我們的父親說：『你們再去給我買些糧來。』
GEN|44|26|我們說：『我們不能下去。最小的弟弟若和我們同去，我們就可以下去。因為，最小的弟弟若不和我們同去，我們必不能見那人的面。』
GEN|44|27|你僕人，我父親對我們說：『你們知道我的妻子給我生了兩個兒子。
GEN|44|28|一個離開我走了，我說他必是被野獸撕碎了，直到如今我再沒有見過他；
GEN|44|29|現在你們又要把這個從我面前帶走。倘若他遭難，那麼你們就害我白髮蒼蒼、悲悲慘慘下陰間去了。』
GEN|44|30|如今我回到你僕人，我父親那裏，若沒有這年輕人和我們同去，我父親的命是與這年輕人的命相連的，
GEN|44|31|當我們的父親看見沒有了這年輕人，他就會死。這樣，我們就害你僕人，我們的父親白髮蒼蒼、悲悲慘慘下陰間去了。
GEN|44|32|僕人曾向我父親為這年輕人擔保，說：『我若不帶他回來交給父親，我就在父親面前永遠擔當這罪。』
GEN|44|33|現在，求你把僕人留下，代替這年輕人作我主的奴隸，讓這年輕人和他哥哥們一同上去。
GEN|44|34|若這年輕人不和我一起，我怎能上到我父親那裏呢？恐怕我要看到災禍臨到我父親了。」
GEN|45|1|約瑟 在所有侍立在他旁邊的人面前情不自禁，就喊叫說：「每一個人都離開我，出去吧！」 約瑟 和兄弟相認的時候沒有一人站在他那裏。
GEN|45|2|他放聲大哭， 埃及 人聽見了，法老家中的人也聽見了。
GEN|45|3|約瑟 對他兄弟們說：「我就是 約瑟 。我的父親還在嗎？」他兄弟們不敢回答他，因為他們在他面前都很驚惶。
GEN|45|4|約瑟 又對他兄弟們說：「靠近我一點。」他們就近前來。他說：「我是被你們賣到 埃及 的兄弟 約瑟 。
GEN|45|5|現在，不要因為把我賣到這裏而憂傷，對自己生氣，因為上帝差我在你們以先來，為要保全性命。
GEN|45|6|現在這地的饑荒已經二年了，還有五年不能耕種，沒有收成。
GEN|45|7|上帝差我在你們以先來，為要給你們在世上存留餘種，大施拯救，保全你們的性命。
GEN|45|8|這樣看來，差我到這裏來的不是你們，而是上帝。他又使我如同法老之父，作他全家之主，和 埃及 全地掌權的人。
GEN|45|9|你們要趕緊上到我父親那裏，對他說：『你兒子 約瑟 這樣說：上帝已立我作全 埃及 之主，請你下到我這裏來，不要耽擱。
GEN|45|10|你和你的兒子孫子，羊群牛群，以及一切所有的，都可以住在 歌珊 地，與我相近。
GEN|45|11|我要在那裏奉養你，因為還有五年的饑荒，免得你和你的家屬，以及一切所有的，都陷入窮困中。』
GEN|45|12|看哪，你們的眼睛和我弟弟 便雅憫 的眼睛都看見，是我親口對你們說話。
GEN|45|13|你們要把我在 埃及 一切的尊榮和你們所有看見的事情都告訴我父親，也要趕緊請我父親下到這裏來。」
GEN|45|14|於是 約瑟 伏在他弟弟 便雅憫 的頸項上哭， 便雅憫 也在他的頸項上哭。
GEN|45|15|他又親眾兄弟，伏著他們哭。過後，他的兄弟就和他說話。
GEN|45|16|這消息傳到法老的宮裏，說：「 約瑟 的兄弟們來了。」法老和他的臣僕眼中都看為好。
GEN|45|17|法老對 約瑟 說：「你要吩咐你的兄弟們說：『你們要這樣做：把馱子抬在牲口上，動身到 迦南 地去，
GEN|45|18|請你們的父親和你們的家屬都到我這裏來，我要把 埃及 地的美物賜給你們，你們也要吃這地肥美的出產。』
GEN|45|19|你要吩咐他們：『要這樣做：從 埃及 地帶著車輛去，把你們的孩子和妻子，以及你們的父親都接來。
GEN|45|20|你們的眼不要顧惜你們的家具，因為 埃及 全地的美物都是你們的。』」
GEN|45|21|以色列 的兒子們就照樣做了。 約瑟 遵照法老的吩咐，給他們車輛和路上需用的食物。
GEN|45|22|他又給所有哥哥每人一套衣服， 卻給 便雅憫 三百銀子，五套衣服。
GEN|45|23|他也送給父親十匹公驢，馱著 埃及 的美物，以及十匹母驢，馱著給他父親在路上需用的穀物、餅和糧食。
GEN|45|24|於是 約瑟 送他的兄弟們回去，對他們說：「你們不要在路上爭吵。」
GEN|45|25|他們從 埃及 上去，來到 迦南 地他們的父親 雅各 那裏，
GEN|45|26|告訴他說：「 約瑟 還活著，並且作了 埃及 全地掌權的人。」 雅各 心裏冰涼，因為不信他們。
GEN|45|27|他們就把 約瑟 對他們所說一切的話都告訴了他。他看見 約瑟 派來接他的車輛，他們父親 雅各 的靈就甦醒了。
GEN|45|28|以色列 說：「夠了！我的兒子 約瑟 還活著，我要趁我未死之前去見他。」
GEN|46|1|以色列 帶著一切所有的，起程到 別是巴 去，獻祭給他父親 以撒 的上帝。
GEN|46|2|夜間，上帝在異象中對 以色列 說：「 雅各 ！ 雅各 ！」他說：「我在這裏。」
GEN|46|3|上帝說：「我是上帝，你父親的上帝。不要害怕下 埃及 去，因為我必使你在那裏成為大國。
GEN|46|4|我要和你同下 埃及 去，也必定帶你上來； 約瑟 要親手合上你的眼睛。」
GEN|46|5|雅各 就從 別是巴 起行。 以色列 的兒子讓他們的父親 雅各 和他們的孩子、妻子都坐在法老為 雅各 派來的車上。
GEN|46|6|他們也帶著 迦南 地所得的牲畜和財物來到 埃及 。 雅各 和他所有的子孫都一同來了。
GEN|46|7|他把他的兒子、孫子、女兒、孫女，他所有的子孫一同帶到 埃及 。
GEN|46|8|這些是來到 埃及 的 以色列 人， 雅各 和他子孫的名字： 雅各 的長子是 呂便 。
GEN|46|9|呂便 的兒子是 哈諾 、 法路 、 希斯倫 、 迦米 。
GEN|46|10|西緬 的兒子是 耶母利 、 雅憫 、 阿轄 、 雅斤 、 瑣轄 ，還有 迦南 女子生的兒子 掃羅 。
GEN|46|11|利未 的兒子是 革順 、 哥轄 、 米拉利 。
GEN|46|12|猶大 的兒子是 珥 、 俄南 、 示拉 、 法勒斯 、 謝拉 ； 珥 與 俄南 死在 迦南 地。 法勒斯 的兒子是 希斯崙 、 哈母勒 。
GEN|46|13|以薩迦 的兒子是 陀拉 、 普瓦 、 約伯 、 伸崙 。
GEN|46|14|西布倫 的兒子是 西烈 、 以倫 、 雅利 。
GEN|46|15|這是 利亞 在 巴旦‧亞蘭 為 雅各 所生的兒孫，還有女兒 底拿 ，兒孫共三十三人。
GEN|46|16|迦得 的兒子是 洗非芸 、 哈基 、 書尼 、 以斯本 、 以利 、 亞羅底 、 亞列利 。
GEN|46|17|亞設 的兒子是 音拿 、 亦施瓦 、 亦施韋 、 比利亞 ，還有他們的妹妹 西拉 。 比利亞 的兒子是 希別 、 瑪結 。
GEN|46|18|這是 拉班 給他女兒 利亞 的婢女 悉帕 的兒孫，她為 雅各 所生的共有十六人。
GEN|46|19|雅各 之妻 拉結 的兒子是 約瑟 和 便雅憫 。
GEN|46|20|約瑟 在 埃及 地生了 瑪拿西 和 以法蓮 ，是 安城 的祭司 波提非拉 的女兒 亞西納 為 約瑟 生的。
GEN|46|21|便雅憫 的兒子是 比拉 、 比結 、 亞實別 、 基拉 、 乃幔 、 以希 、 羅實 、 母平 、 戶平 、 亞勒 。
GEN|46|22|這是 拉結 為 雅各 所生的兒孫，共有十四人。
GEN|46|23|但 的兒子是 戶伸 。
GEN|46|24|拿弗他利 的兒子是 雅薛 、 沽尼 、 耶色 、 示冷 。
GEN|46|25|這是 拉班 給他女兒 拉結 的婢女 辟拉 的兒孫，她為 雅各 所生的共有七人。
GEN|46|26|那與 雅各 同到 埃及 的，除了他媳婦之外，凡從他生的共有六十六人。
GEN|46|27|還有 約瑟 在 埃及 所生的兩個兒子。到 埃及 的 雅各 全家共有七十人。
GEN|46|28|雅各 派 猶大 先到 約瑟 那裏，請他先指示到 歌珊 去的路；於是他們來到了 歌珊 地。
GEN|46|29|約瑟 備好座車，上 歌珊 去迎接他的父親 以色列 。他見到父親，就伏在父親的頸項上，在父親的頸項上哭了許久。
GEN|46|30|以色列 對 約瑟 說：「我見了你的面，知道你還活著，現在我可以死了。」
GEN|46|31|約瑟 對他兄弟和他父親的全家說：「我要上去告訴法老，對他說：『我在 迦南 地的兄弟和我父親的全家，都到我這裏來了。
GEN|46|32|他們是牧羊人，是牧放牲畜的人；他們把羊群牛群和一切所有的都帶來了。』
GEN|46|33|等到法老召見你們，說：『你們是做甚麼的？』
GEN|46|34|你們就說：『你的僕人，從幼年直到現在，都是牧放牲畜的人，我們和我們的祖宗都是這樣。』如此，你們就可以住在 歌珊 地，因為凡牧羊的都被 埃及 人厭惡。」
GEN|47|1|約瑟 進去告訴法老說：「我的父親和我的兄弟帶著羊群牛群，以及他們一切所有的，從 迦南 地來了。看哪，他們正在 歌珊 地。」
GEN|47|2|約瑟 從他所有兄弟中挑選五個人，引他們到法老面前。
GEN|47|3|法老對 約瑟 的兄弟說：「你們是做甚麼的？」他們對法老說：「你僕人是牧羊的，我們和我們的祖宗都是這樣。」
GEN|47|4|他們又對法老說：「 迦南 地的饑荒非常嚴重，僕人的羊群沒有牧草，所以我們來到這地寄居。現在求你准許僕人住在 歌珊 地。」
GEN|47|5|法老對 約瑟 說：「你的父親和你的兄弟到你這裏來了，
GEN|47|6|埃及 地都在你面前，只管讓你父親和你兄弟住在最好的地，他們可以住在 歌珊 地。你若知道他們中間有能幹的人，就派他們看管我的牲畜。」
GEN|47|7|約瑟 帶他父親 雅各 來，站在法老面前， 雅各 就為法老祝福。
GEN|47|8|法老對 雅各 說：「你平生的年日是多少呢？」
GEN|47|9|雅各 對法老說：「我在世寄居的年日是一百三十年，我一生的歲月又短又苦，比不上我祖先在世寄居的年日。」
GEN|47|10|雅各 又為法老祝福，就從法老面前退出去了。
GEN|47|11|約瑟 安頓他的父親和兄弟，遵照法老的命令，把 埃及 境內最好的地，就是 蘭塞 地，給他們作為產業。
GEN|47|12|約瑟 用糧食供給他父親和兄弟們，以及他父親全家的人，照扶養親屬的人口供給。
GEN|47|13|饑荒非常嚴重，全地都絕了糧， 埃及 地和 迦南 地都因饑荒耗損了。
GEN|47|14|約瑟 收集了 埃及 地和 迦南 地所有的銀子，就是眾人買糧的銀子， 約瑟 就把那些銀子都帶到法老的宮裏。
GEN|47|15|埃及 地和 迦南 地的銀子都花光了， 埃及 眾人到 約瑟 那裏，說：「我們的銀子都用完了，求你給我們糧食吧！我們為甚麼要死在你面前呢？」
GEN|47|16|約瑟 說：「銀子若是用完了，可以把你們的牲畜賣給我，我就以你們的牲畜換糧食給你們。」
GEN|47|17|於是他們把牲畜帶到 約瑟 那裏， 約瑟 就拿糧食換了他們的馬、羊、牛、驢；那一年他因換他們一切的牲畜，用糧食養活他們。
GEN|47|18|那一年過去，第二年他們又來到 約瑟 那裏，對他說：「不瞞我主，我們的銀子都花光了，牲畜也都歸於我主了。我們在我主面前，除了自己的身體和土地以外，一無所剩。
GEN|47|19|你為甚麼要眼看著我們人死地荒呢？求你用糧食買我們和我們的地，我們和我們的地就要為法老效力。求你給我們種子，使我們可以存活，不致死亡，土地也不致荒蕪。」
GEN|47|20|於是， 約瑟 為法老買了 埃及 所有的土地， 埃及 人因饑荒所迫，都賣了自己的田地；那些地都歸給法老了。
GEN|47|21|至於百姓，從 埃及 邊界的一端到另一端， 約瑟 使他們作奴隸。
GEN|47|22|只有祭司的土地， 約瑟 沒有買，因為祭司從法老領取薪俸，靠法老的薪俸過活，所以沒有賣自己的土地。
GEN|47|23|約瑟 對百姓說：「看哪，我今日為法老買了你們和你們的土地。看，這些種子是給你們的，你們可以耕種土地。
GEN|47|24|將來收割的時候，你們要把五分之一納給法老，另外四分可以給你們作田地的種子，作你們和你們全家大小的食物。」
GEN|47|25|他們說：「你救了我們的性命，願我們在我主眼前蒙恩，我們情願作法老的奴隸。」
GEN|47|26|於是 約瑟 為 埃及 的土地立下定例，直到今日，就是收成的五分之一要歸法老。惟獨祭司的土地例外，不歸於法老。
GEN|47|27|以色列 人住在 埃及 境內的 歌珊 地。他們在那裏得了產業，並且生養眾多。
GEN|47|28|雅各 住在 埃及 地十七年。 雅各 一生的年日是一百四十七年。
GEN|47|29|以色列 的死期快到了，就叫了他兒子 約瑟 來，對他說：「我若在你眼前蒙恩，把你的手放在我大腿底下，以慈愛和誠實向我承諾，必不將我葬在 埃及 。
GEN|47|30|我與我祖先同睡的時候，你要將我帶出 埃及 ，把我葬在他們所葬的地方。」 約瑟 說：「我必遵照你的吩咐去做。」
GEN|47|31|雅各 說：「你向我起誓吧！」 約瑟 就向他起了誓。於是 以色列 在床頭 敬拜。
GEN|48|1|這些事以後，有人告訴 約瑟 說：「看哪，你的父親病了。」他就帶著兩個兒子 瑪拿西 和 以法蓮 同去。
GEN|48|2|有人告訴 雅各 說：「看哪，你的兒子 約瑟 到你這裏來了。」 以色列 就勉強在床上坐起來。
GEN|48|3|雅各 對 約瑟 說：「全能的上帝曾在 迦南 地的 路斯 向我顯現，賜福給我，
GEN|48|4|對我說：『看哪，我必使你生養眾多，成為許多民族，又要將這地賜給你的後裔，永遠為業。』
GEN|48|5|我未到 埃及 你那裏之前，你在 埃及 地所生的 以法蓮 和 瑪拿西 這兩個兒子，現在他們是我的，正如 呂便 和 西緬 是我的一樣。
GEN|48|6|你在他們以後所生的後裔就是你的，這些後裔可以在自己兄弟的名下得產業。
GEN|48|7|至於我，我從 巴旦 回來的時候， 拉結 在我身旁死了，就是在往 迦南 地的路上，離 以法他 還有一段路程。我就把她葬在往 以法他 的路旁； 以法他 就是 伯利恆 。」
GEN|48|8|以色列 看見 約瑟 的兒子，就說：「這些是誰？」
GEN|48|9|約瑟 對他父親說：「這是上帝在這裏賜給我的兒子。」 以色列 說：「領他們到我跟前，我要為他們祝福。」
GEN|48|10|以色列 年紀老邁，眼睛昏花，不能看見。 約瑟 領他們到他跟前，他就和他們親吻，抱著他們。
GEN|48|11|以色列 對 約瑟 說：「我沒有想到能夠見你的面。看哪，上帝還讓我看見你的兒子。」
GEN|48|12|約瑟 把他們從 以色列 兩膝中間領出來，自己臉伏於地下拜。
GEN|48|13|然後， 約瑟 牽著他們兩個，帶到父親跟前，右手牽 以法蓮 到 以色列 的左邊，左手牽 瑪拿西 到 以色列 的右邊。
GEN|48|14|以色列 卻伸出右手來，按在次子 以法蓮 的頭上，又交叉伸出左手來，按在長子 瑪拿西 的頭上。
GEN|48|15|他就為 約瑟 祝福說： 「願我祖父 亞伯拉罕 和我父親 以撒 所事奉的上帝， 就是一生牧養我直到今日的上帝，
GEN|48|16|救贖我脫離一切患難的那位使者，賜福給這兩個孩子。 願我的名，我祖父 亞伯拉罕 和我父親 以撒 的名藉著他們得以流傳。 又願他們在全地上多多繁衍。」
GEN|48|17|約瑟 見父親把右手按在 以法蓮 的頭上，他看為不好，就提起他父親的手，要從 以法蓮 的頭上移到 瑪拿西 的頭上。
GEN|48|18|約瑟 對父親說：「我父，不是這樣。這個才是長子，請你把右手按在他頭上。」
GEN|48|19|他父親卻不肯，說：「我知道，我兒，我知道。他也要成為一族，也要強大。可是他的弟弟將來比他還要強大；他弟弟的後裔要成為許多國家。」
GEN|48|20|以色列 就在當日為他們祝福，說：「 以色列 人要指著你們祝福，說：『願上帝使你如 以法蓮 、 瑪拿西 一樣。』」於是他立 以法蓮 在 瑪拿西 之上。
GEN|48|21|以色列 又對 約瑟 說：「看哪，我快要死了，但上帝必與你們同在，領你們回到你們祖先之地。
GEN|48|22|從前我用刀用弓從 亞摩利 人手下奪取的那一份，我要把它賜給你，使你比你的兄弟多得一份 。」
GEN|49|1|雅各 叫了他的兒子來，說：「你們都來聚集，讓我把你們日後要遇到的事告訴你們。
GEN|49|2|雅各 的兒子們，你們要聚集，要聆聽， 聽你們父親 以色列 的話。
GEN|49|3|呂便 啊，你是我的長子，我的力量， 我壯年頭生之子， 極有尊榮，權力超群。
GEN|49|4|你卻放縱如水，必不得居首位； 因為你上了你父親的床， 你 上了我的榻，污辱了它！
GEN|49|5|西緬 和 利未 是兄弟； 他們的刀劍是殘暴的兵器。
GEN|49|6|願我的心不與他們同謀， 願我的靈 不與他們合夥； 因為他們在烈怒中殺人， 任意割斷牛腿的筋。
GEN|49|7|他們火爆的烈怒可詛， 他們兇殘的憤恨可咒！ 我要把他們分散在 雅各 中， 使他們散居在 以色列 。
GEN|49|8|猶大 啊，你的兄弟必讚美你， 你的手必掐住仇敵的頸項， 你父親的兒子要向你下拜。
GEN|49|9|猶大 是隻小獅子； 我兒啊，你捕獲了獵物就上去。 他蹲伏，他躺臥，如公獅， 又如母獅，誰敢惹他呢？
GEN|49|10|權杖必不離 猶大 ， 統治者的杖必不離他兩腳之間， 直等細羅 來到， 萬民都要歸順他。
GEN|49|11|猶大 把小驢拴在葡萄樹上， 把驢駒拴在佳美的葡萄樹上。 他在葡萄酒中洗衣服， 在葡萄汁 中洗長袍。
GEN|49|12|他的眼睛比 酒紅潤， 他的牙齒比奶潔白。
GEN|49|13|西布倫 必住在海邊， 必成為停船的港口； 他的疆界必延到 西頓 。
GEN|49|14|以薩迦 是匹強壯的驢， 臥在羊圈之中。
GEN|49|15|他看見居所安舒， 土地肥美， 就屈肩負重， 成為服勞役的僕人。
GEN|49|16|但 必為他的百姓伸冤 ， 作為 以色列 支派之一。
GEN|49|17|但 必作道旁的蛇， 路邊的毒蛇， 咬傷馬蹄， 使騎馬的人向後墜落。
GEN|49|18|耶和華啊，我等候你的救恩。
GEN|49|19|迦得 必被襲擊者襲擊 ， 他卻要襲擊他們的腳跟。
GEN|49|20|亞設 必出豐盛的糧食， 要供應君王的佳肴。
GEN|49|21|拿弗他利 是被釋放的母鹿， 他要生出可愛的小鹿 。
GEN|49|22|約瑟 是多結果子的樹枝， 是泉旁多結果的枝子； 他的枝條伸出牆外。
GEN|49|23|弓箭手惡意攻擊他， 敵對他，向他射箭。
GEN|49|24|但他的弓仍舊堅硬， 他的手臂靈活敏捷， 這是因 雅各 的大能者的手， 從那裏，他是 以色列 的牧者， 以色列 的磐石 。
GEN|49|25|你父親的上帝必幫助你； 全能者必賜福給你： 天上的福， 深淵下面蘊藏的福， 以及生育哺養的福。
GEN|49|26|你父親的福 勝過我祖先的福， 直到永世山嶺的極限。 這些福必降在 約瑟 的頭上， 臨到那與兄弟有分別之人的頭頂上。
GEN|49|27|便雅憫 是隻抓撕掠物的狼， 早晨要吃他的獵物， 晚上要分他的擄物。」
GEN|49|28|這一切是 以色列 的十二個支派。這是他們的父親對他們所說的話，他按照各人的福分為他們祝福。
GEN|49|29|他又吩咐他們說：「我快要歸到我祖先 那裏。你們要將我葬在 赫 人 以弗崙 田間的洞裏，與我的祖先在一處，
GEN|49|30|就是在 迦南 地 幔利 對面的 麥比拉 田間的洞裏，那田是 亞伯拉罕 向 赫 人 以弗崙 買來作墳地的產業。
GEN|49|31|亞伯拉罕 和他的妻子 撒拉 葬在那裏； 以撒 和他的妻子 利百加 也葬在那裏。我也在那裏葬了 利亞 。
GEN|49|32|那塊田和田間的洞是向 赫 人買的。」
GEN|49|33|雅各 囑咐眾子完畢後，就把腳收在床上斷了氣，歸到他祖先 那裏去了。
GEN|50|1|約瑟 伏在他父親的臉上，在他臉上哭，又親他。
GEN|50|2|約瑟 吩咐伺候他的醫生們用香料塗他父親，醫生就用香料塗了 以色列 。
GEN|50|3|四十天滿了，就是塗香料所規定的日子滿了。 埃及 人為他哀哭了七十天。
GEN|50|4|過了哀悼的日子， 約瑟 對法老家中的人說：「我若在你們眼前蒙恩，請你們對法老說：
GEN|50|5|『我父親曾叫我起誓說：看哪，我快要死了，你要將我葬在 迦南 地，在我為自己所掘的墳墓裏。』現在求你准我上去葬我父親，然後我必回來。」
GEN|50|6|法老說：「你可以上去，照你父親叫你起的誓，將他安葬。」
GEN|50|7|於是 約瑟 上去葬他父親。與他一同上去的有法老的眾臣僕和法老家中的長老，以及 埃及 地所有的長老，
GEN|50|8|還有 約瑟 的全家和他的兄弟們，以及他父親的家屬；只留下他們的孩子和羊群牛群在 歌珊 地。
GEN|50|9|又有車輛和駕駛兵和他一同上去，隊伍非常龐大。
GEN|50|10|他們到了 約旦河 東 亞達 的禾場，就在那裏大大地號咷痛哭。 約瑟 為他父親哀哭了七天。
GEN|50|11|迦南 的居民看見 亞達 禾場上的哀哭，就說：「這是 埃及 人一場極大的哀哭。」因此那地方名叫 亞伯‧麥西 ，是在 約旦河 東。
GEN|50|12|雅各 的兒子們遵照父親的吩咐去辦了，
GEN|50|13|他們把他送到 迦南 地，葬在 幔利 對面的 麥比拉 田間的洞裏；那田是 亞伯拉罕 向 赫 人 以弗崙 買來作墳地的產業。
GEN|50|14|約瑟 葬了他父親以後，就和他的兄弟，以及所有同他上去葬他父親的人，都回 埃及 去了。
GEN|50|15|約瑟 的哥哥們見父親死了，就說：「也許 約瑟 仍然懷恨我們，會照我們從前待他一切的惡，重重報復我們。」
GEN|50|16|他們就傳口信給 約瑟 說：「你父親未死之前曾吩咐說：
GEN|50|17|『你們要對 約瑟 這樣說：從前你哥哥們惡待你，你要饒恕他們的過犯和罪惡。』現在求你饒恕你父親的上帝之僕人們的過犯。」他們對 約瑟 說了這話， 約瑟 就哭了。
GEN|50|18|他的哥哥們又來俯伏在他面前，說：「看哪，我們是你的奴隸。」
GEN|50|19|約瑟 對他們說：「不要怕，我豈能代替上帝呢？
GEN|50|20|從前你們的意思是要害我，但上帝的意思原是好的，要使許多百姓得以存活，成就今日的光景。
GEN|50|21|現在你們不要害怕，我必養活你們和你們的孩子。」於是 約瑟 安慰他們，講了使他們安心的話。
GEN|50|22|約瑟 和他父親的家屬都住在 埃及 。 約瑟 活了一百一十年。
GEN|50|23|約瑟 看到 以法蓮 第三代的子孫。 瑪拿西 的孫子， 瑪吉 的兒子，出生時都放在 約瑟 的膝上。
GEN|50|24|約瑟 對他的兄弟說：「我快要死了，但上帝必定看顧你們，領你們從這地上去，到他起誓應許給 亞伯拉罕 、 以撒 、 雅各 之地。」
GEN|50|25|約瑟 叫 以色列 的子孫起誓：「上帝必定眷顧你們，你們要把我的骸骨從這裏帶上去。」
GEN|50|26|約瑟 死了，那時他一百一十歲。人用香料塗了他，把他收殮在棺材裏，停放在 埃及 。
