LAM|1|1|How lonely sits the citythat was full of people! How like a widow has she become, she who was great among the nations! She who was a princess among the provinces has become a slave.
LAM|1|2|She weeps bitterly in the night, with tears on her cheeks; among all her lovers she has none to comfort her; all her friends have dealt treacherously with her; they have become her enemies.
LAM|1|3|Judah has gone into exile because of affliction and hard servitude; she dwells now among the nations, but finds no resting place; her pursuers have all overtaken her in the midst of her distress.
LAM|1|4|The roads to Zion mourn, for none come to the festival; all her gates are desolate; her priests groan; her virgins have been afflicted, and she herself suffers bitterly.
LAM|1|5|Her foes have become the head; her enemies prosper, because the LORD has afflicted her for the multitude of her transgressions; her children have gone away, captives before the foe.
LAM|1|6|From the daughter of Zion all her majesty has departed. Her princes have become like deer that find no pasture; they fled without strength before the pursuer.
LAM|1|7|Jerusalem remembers in the days of her affliction and wandering all the precious things that were hers from days of old. When her people fell into the hand of the foe, and there was none to help her, her foes gloated over her; they mocked at her downfall.
LAM|1|8|Jerusalem sinned grievously; therefore she became filthy; all who honored her despise her, for they have seen her nakedness; she herself groans and turns her face away.
LAM|1|9|Her uncleanness was in her skirts; she took no thought of her future; therefore her fall is terrible; she has no comforter. "O LORD, behold my affliction, for the enemy has triumphed!"
LAM|1|10|The enemy has stretched out his hands over all her precious things; for she has seen the nations enter her sanctuary, those whom you forbade to enter your congregation.
LAM|1|11|All her people groan as they search for bread; they trade their treasures for food to revive their strength. "Look, O LORD, and see, for I am despised."
LAM|1|12|"Is it nothing to you, all you who pass by? Look and see if there is any sorrow like my sorrow, which was brought upon me, which the LORD inflicted on the day of his fierce anger.
LAM|1|13|"From on high he sent fire; into my bones he made it descend; he spread a net for my feet; he turned me back; he has left me stunned, faint all the day long.
LAM|1|14|"My transgressions were bound into a yoke; by his hand they were fastened together; they were set upon my neck; he caused my strength to fail; the Lord gave me into the hands of those whom I cannot withstand.
LAM|1|15|"The Lord rejected all my mighty men in my midst; he summoned an assembly against me to crush my young men; the Lord has trodden as in a winepress the virgin daughter of Judah.
LAM|1|16|"For these things I weep; my eyes flow with tears; for a comforter is far from me, one to revive my spirit; my children are desolate, for the enemy has prevailed."
LAM|1|17|Zion stretches out her hands, but there is none to comfort her; the LORD has commanded against Jacob that his neighbors should be his foes; Jerusalem has become a filthy thing among them.
LAM|1|18|"The LORD is in the right, for I have rebelled against his word; but hear, all you peoples, and see my suffering; my young women and my young men have gone into captivity.
LAM|1|19|"I called to my lovers, but they deceived me; my priests and elders perished in the city, while they sought food to revive their strength.
LAM|1|20|"Look, O LORD, for I am in distress; my stomach churns; my heart is wrung within me, because I have been very rebellious. In the street the sword bereaves; in the house it is like death.
LAM|1|21|"They heard my groaning, yet there is no one to comfort me. All my enemies have heard of my trouble; they are glad that you have done it. You have brought the day you announced; now let them be as I am.
LAM|1|22|"Let all their evildoing come before you, and deal with them as you have dealt with me because of all my transgressions; for my groans are many, and my heart is faint."
LAM|2|1|How the Lord in his anger has set the daughter of Zion under a cloud! He has cast down from heaven to earth the splendor of Israel; he has not remembered his footstool in the day of his anger.
LAM|2|2|The Lord has swallowed up without mercy all the habitations of Jacob; in his wrath he has broken down the strongholds of the daughter of Judah; he has brought down to the ground in dishonor the kingdom and its rulers.
LAM|2|3|He has cut down in fierce anger all the might of Israel; he has withdrawn from them his right hand in the face of the enemy; he has burned like a flaming fire in Jacob, consuming all around.
LAM|2|4|He has bent his bow like an enemy, with his right hand set like a foe; and he has killed all who were delightful in our eyes in the tent of the daughter of Zion; he has poured out his fury like fire.
LAM|2|5|The Lord has become like an enemy; he has swallowed up Israel; he has swallowed up all its palaces; he has laid in ruins its strongholds, and he has multiplied in the daughter of Judah mourning and lamentation.
LAM|2|6|He has laid waste his booth like a garden, laid in ruins his meeting place; the LORD has made Zion forget festival and Sabbath, and in his fierce indignation has spurned king and priest.
LAM|2|7|The Lord has scorned his altar, disowned his sanctuary; he has delivered into the hand of the enemy the walls of her palaces; they raised a clamor in the house of the LORD as on the day of festival.
LAM|2|8|The LORD determined to lay in ruins the wall of the daughter of Zion; he stretched out the measuring line; he did not restrain his hand from destroying; he caused rampart and wall to lament; they languished together.
LAM|2|9|Her gates have sunk into the ground; he has ruined and broken her bars; her king and princes are among the nations; the law is no more, and her prophets find no vision from the LORD.
LAM|2|10|The elders of the daughter of Zion sit on the ground in silence; they have thrown dust on their heads and put on sackcloth; the young women of Jerusalem have bowed their heads to the ground.
LAM|2|11|My eyes are spent with weeping; my stomach churns; my bile is poured out to the ground because of the destruction of the daughter of my people, because infants and babies faint in the streets of the city.
LAM|2|12|They cry to their mothers, "Where is bread and wine?" as they faint like a wounded man in the streets of the city, as their life is poured out on their mothers' bosom.
LAM|2|13|What can I say for you, to what compare you, O daughter of Jerusalem? What can I liken to you, that I may comfort you, O virgin daughter of Zion? For your ruin is vast as the sea; who can heal you?
LAM|2|14|Your prophets have seen for you false and deceptive visions; they have not exposed your iniquity to restore your fortunes, but have seen for you oracles that are false and misleading.
LAM|2|15|All who pass along the way clap their hands at you; they hiss and wag their heads at the daughter of Jerusalem; "Is this the city that was called the perfection of beauty, the joy of all the earth?"
LAM|2|16|All your enemies rail against you; they hiss, they gnash their teeth, they cry: "We have swallowed her! Ah, this is the day we longed for; now we have it; we see it!"
LAM|2|17|The LORD has done what he purposed; he has carried out his word, which he commanded long ago; he has thrown down without pity; he has made the enemy rejoice over you and exalted the might of your foes.
LAM|2|18|Their heart cried to the Lord. O wall of the daughter of Zion, let tears stream down like a torrent day and night! Give yourself no rest, your eyes no respite!
LAM|2|19|"Arise, cry out in the night, at the beginning of the night watches! Pour out your heart like water before the presence of the Lord! Lift your hands to him for the lives of your children, who faint for hunger at the head of every street."
LAM|2|20|Look, O LORD, and see! With whom have you dealt thus? Should women eat the fruit of their womb, the children of their tender care? Should priest and prophet be killed in the sanctuary of the Lord?
LAM|2|21|In the dust of the streets lie the young and the old; my young women and my young men have fallen by the sword; you have killed them in the day of your anger, slaughtering without pity.
LAM|2|22|You summoned as if to a festival day my terrors on every side, and on the day of the anger of the LORD no one escaped or survived; those whom I held and raised my enemy destroyed.
LAM|3|1|I am the man who has seen affliction under the rod of his wrath;
LAM|3|2|he has driven and brought me into darkness without any light;
LAM|3|3|surely against me he turns his hand again and again the whole day long.
LAM|3|4|He has made my flesh and my skin waste away; he has broken my bones;
LAM|3|5|he has besieged and enveloped me with bitterness and tribulation;
LAM|3|6|he has made me dwell in darkness like the dead of long ago.
LAM|3|7|He has walled me about so that I cannot escape; he has made my chains heavy;
LAM|3|8|though I call and cry for help, he shuts out my prayer;
LAM|3|9|he has blocked my ways with blocks of stones; he has made my paths crooked.
LAM|3|10|He is a bear lying in wait for me, a lion in hiding;
LAM|3|11|he turned aside my steps and tore me to pieces; he has made me desolate;
LAM|3|12|he bent his bow and set me as a target for his arrow.
LAM|3|13|He drove into my kidneys the arrows of his quiver;
LAM|3|14|I have become the laughingstock of all peoples, the object of their taunts all day long.
LAM|3|15|He has filled me with bitterness; he has sated me with wormwood.
LAM|3|16|He has made my teeth grind on gravel, and made me cower in ashes;
LAM|3|17|my soul is bereft of peace; I have forgotten what happiness is;
LAM|3|18|so I say, "My endurance has perished; so has my hope from the LORD."
LAM|3|19|Remember my affliction and my wanderings, the wormwood and the gall!
LAM|3|20|My soul continually remembers it and is bowed down within me.
LAM|3|21|But this I call to mind, and therefore I have hope:
LAM|3|22|The steadfast love of the LORD never ceases; his mercies never come to an end;
LAM|3|23|they are new every morning; great is your faithfulness.
LAM|3|24|"The LORD is my portion," says my soul, "therefore I will hope in him."
LAM|3|25|The LORD is good to those who wait for him, to the soul who seeks him.
LAM|3|26|It is good that one should wait quietly for the salvation of the LORD.
LAM|3|27|It is good for a man that he bear the yoke in his youth.
LAM|3|28|Let him sit alone in silence when it is laid on him;
LAM|3|29|let him put his mouth in the dust- there may yet be hope;
LAM|3|30|let him give his cheek to the one who strikes, and let him be filled with insults.
LAM|3|31|For the Lord will not cast off forever,
LAM|3|32|but, though he cause grief, he will have compassion according to the abundance of his steadfast love;
LAM|3|33|for he does not willingly afflict or grieve the children of men.
LAM|3|34|To crush underfoot all the prisoners of the earth,
LAM|3|35|to deny a man justice in the presence of the Most High,
LAM|3|36|to subvert a man in his lawsuit, the Lord does not approve.
LAM|3|37|Who has spoken and it came to pass, unless the Lord has commanded it?
LAM|3|38|Is it not from the mouth of the Most High that good and bad come?
LAM|3|39|Why should a living man complain, a man, about the punishment of his sins?
LAM|3|40|Let us test and examine our ways, and return to the LORD!
LAM|3|41|Let us lift up our hearts and hands to God in heaven:
LAM|3|42|"We have transgressed and rebelled, and you have not forgiven.
LAM|3|43|"You have wrapped yourself with anger and pursued us, killing without pity;
LAM|3|44|you have wrapped yourself with a cloud so that no prayer can pass through.
LAM|3|45|You have made us scum and garbage among the peoples.
LAM|3|46|"All our enemies open their mouths against us;
LAM|3|47|panic and pitfall have come upon us, devastation and destruction;
LAM|3|48|my eyes flow with rivers of tears because of the destruction of the daughter of my people.
LAM|3|49|"My eyes will flow without ceasing, without respite,
LAM|3|50|until the LORD from heaven looks down and sees;
LAM|3|51|my eyes cause me grief at the fate of all the daughters of my city.
LAM|3|52|"I have been hunted like a bird by those who were my enemies without cause;
LAM|3|53|they flung me alive into the pit and cast stones on me;
LAM|3|54|water closed over my head; I said, 'I am lost.'
LAM|3|55|"I called on your name, O LORD, from the depths of the pit;
LAM|3|56|you heard my plea, 'Do not close your ear to my cry for help!'
LAM|3|57|You came near when I called on you; you said, 'Do not fear!'
LAM|3|58|"You have taken up my cause, O Lord; you have redeemed my life.
LAM|3|59|You have seen the wrong done to me, O LORD; judge my cause.
LAM|3|60|You have seen all their vengeance, all their plots against me.
LAM|3|61|"You have heard their taunts, O LORD, all their plots against me.
LAM|3|62|The lips and thoughts of my assailants are against me all the day long.
LAM|3|63|Behold their sitting and their rising; I am the object of their taunts.
LAM|3|64|"You will repay them, O LORD, according to the work of their hands.
LAM|3|65|You will give them dullness of heart; your curse will be on them.
LAM|3|66|You will pursue them in anger and destroy them from under your heavens, O LORD."
LAM|4|1|How the gold has grown dim, how the pure gold is changed! The holy stones lie scattered at the head of every street.
LAM|4|2|The precious sons of Zion, worth their weight in fine gold, how they are regarded as earthen pots, the work of a potter's hands!
LAM|4|3|Even jackals offer the breast; they nurse their young, but the daughter of my people has become cruel, like the ostriches in the wilderness.
LAM|4|4|The tongue of the nursing infant sticks to the roof of its mouth for thirst; the children beg for food, but no one gives to them.
LAM|4|5|Those who once feasted on delicacies perish in the streets; those who were brought up in purple embrace ash heaps.
LAM|4|6|For the chastisement of the daughter of my people has been greater than the punishment of Sodom, which was overthrown in a moment, and no hands were wrung for her.
LAM|4|7|Her princes were purer than snow, whiter than milk; their bodies were more ruddy than coral, the beauty of their form was like sapphire.
LAM|4|8|Now their face is blacker than soot; they are not recognized in the streets; their skin has shriveled on their bones; it has become as dry as wood.
LAM|4|9|Happier were the victims of the sword than the victims of hunger, who wasted away, pierced by lack of the fruits of the field.
LAM|4|10|The hands of compassionate women have boiled their own children; they became their food during the destruction of the daughter of my people.
LAM|4|11|The LORD gave full vent to his wrath; he poured out his hot anger, and he kindled a fire in Zion that consumed its foundations.
LAM|4|12|The kings of the earth did not believe, nor any of the inhabitants of the world, that foe or enemy could enter the gates of Jerusalem.
LAM|4|13|This was for the sins of her prophets and the iniquities of her priests, who shed in the midst of her the blood of the righteous.
LAM|4|14|They wandered, blind, through the streets; they were so defiled with blood that no one was able to touch their garments.
LAM|4|15|"Away! Unclean!" people cried at them. "Away! Away! Do not touch!" So they became fugitives and wanderers; people said among the nations, "They shall stay with us no longer."
LAM|4|16|The LORD himself has scattered them; he will regard them no more; no honor was shown to the priests, no favor to the elders.
LAM|4|17|Our eyes failed, ever watching vainly for help; in our watching we watched for a nation which could not save.
LAM|4|18|They dogged our steps so that we could not walk in our streets; our end drew near; our days were numbered, for our end had come.
LAM|4|19|Our pursuers were swifter than the eagles in the heavens; they chased us on the mountains; they lay in wait for us in the wilderness.
LAM|4|20|The breath of our nostrils, the LORD's anointed, was captured in their pits, of whom we said, "Under his shadow we shall live among the nations."
LAM|4|21|Rejoice and be glad, O daughter of Edom, you who dwell in the land of Uz; but to you also the cup shall pass; you shall become drunk and strip yourself bare.
LAM|4|22|The punishment of your iniquity, O daughter of Zion, is accomplished; he will keep you in exile no longer; but your iniquity, O daughter of Edom, he will punish; he will uncover your sins.
LAM|5|1|Remember, O LORD, what has befallen us; look, and see our disgrace!
LAM|5|2|Our inheritance has been turned over to strangers, our homes to foreigners.
LAM|5|3|We have become orphans, fatherless; our mothers are like widows.
LAM|5|4|We must pay for the water we drink; the wood we get must be bought.
LAM|5|5|Our pursuers are at our necks; we are weary; we are given no rest.
LAM|5|6|We have given the hand to Egypt, and to Assyria, to get bread enough.
LAM|5|7|Our fathers sinned, and are no more; and we bear their iniquities.
LAM|5|8|Slaves rule over us; there is none to deliver us from their hand.
LAM|5|9|We get our bread at the peril of our lives, because of the sword in the wilderness.
LAM|5|10|Our skin is hot as an oven with the burning heat of famine.
LAM|5|11|Women are raped in Zion, young women in the towns of Judah.
LAM|5|12|Princes are hung up by their hands; no respect is shown to the elders.
LAM|5|13|Young men are compelled to grind at the mill, and boys stagger under loads of wood.
LAM|5|14|The old men have left the city gate, the young men their music.
LAM|5|15|The joy of our hearts has ceased; our dancing has been turned to mourning.
LAM|5|16|The crown has fallen from our head; woe to us, for we have sinned!
LAM|5|17|For this our heart has become sick, for these things our eyes have grown dim,
LAM|5|18|for Mount Zion which lies desolate; jackals prowl over it.
LAM|5|19|But you, O LORD, reign forever; your throne endures to all generations.
LAM|5|20|Why do you forget us forever, why do you forsake us for so many days?
LAM|5|21|Restore us to yourself, O LORD, that we may be restored! Renew our days as of old-
LAM|5|22|unless you have utterly rejected us, and you remain exceedingly angry with us.
